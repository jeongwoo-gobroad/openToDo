                                                                ����  us/       Birthday    @VZ�U   WZ�U  �WZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  pgZ�U  �9����  w/       Workout �U  �m_�U  Pn_�U  �n_Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �r_�U  �g����  ��/      Appointment  �Y�U  ��Y�U  ��YThis_stuffs_This_stuffs_ �U  P�Y�U  �Y�U  ��Y�U  ��Y�U  ������  e�/       Meeting     �sY�U  `tY�U  xYSome_stuffs_Some_stuffs_ �U   �Y�U  ��Y�U  ��Y�U  ��Y�U  �����  ��/       Birthday U  �E[�U  0F[�U  �F[Some_stuffs_Some_stuffs_ �U  �I[�U  pJ[�U  0K[�U  �K[�U  ����  ��/       Birthday    ��\�U  p�\�U  0�\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �\�U  �'����  Z�/      Meeting     �n\�U  @o\�U  �o\Some_stuffs_Some_stuffs_ �U  �r\�U  @s\�U   t\�U  �t\�U  ��S���  e/      Birthday nt ��[�U  0�[�U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p�[�U  ������  �3/       Meeting      �Y�U  ��Y�U  ��YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  $�����  84/      Appointment pmZ�U  0nZ�U  �nZSome_stuffs_Some_stuffs_ �U  p}Z�U  �}Z�U  �rZ�U  psZ�U  @�|���  h_/       Some_stuffs �eY�U  `fY�U  �iYSome_stuffs_Some_stuffs_ �U  �sY�U  `tY�U  xY�U  �xY�U  ����  �/       Appointment @�Z�U  ��Z�U  ��ZThis_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  ��Z�U  X&���  �/       Workout     �[�U  0�[�U  ��[This_stuffs_This_stuffs_ �U  p�[�U  0�[�U  ��[�U  0�[�U  V�&���  ��/      Meeting     �\�U  `\�U   \Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �\�U  �c����  ��/       Meeting     �0Z�U  p1Z�U  02ZSome_stuffs_Some_stuffs_ �U  �4Z�U  0?Z�U  7Z�U  �7Z�U  �w����  ��/      Some_stuffs ��Y�U  p�Y�U  ��YThis_stuffs_This_stuffs_ �U  �Y�U  ��Y�U   �Y�U  �Y�U  �37���  ��/      Appointment �?\�U  �@\�U  @A\Some_stuffs_Some_stuffs_ �U   D\�U  �D\�U  0E\�U  �E\�U  �o����  -�/       Some_stuffs �?Z�U  �@Z�U  PAZThis_stuffs_This_stuffs_ �U  DZ�U  �DZ�U  �EZ�U  PFZ�U  �����  �/      Some_stuffs p@[�U  �@[�U  �A[This_stuffs_This_stuffs_ �U  0D[�U  �D[�U  �E[�U  0F[�U  pGe���  /       Birthday    EY�U  �EY�U  �HYThis_stuffs_This_stuffs_ �U  �PY�U  @QY�U  0TY�U   VY�U  m3����  �&/      Birthday nt  o[�U  �o[�U  @p[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �t[�U  ����  5J/       Appointment �[�U  �[�U   [This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p8[�U  �I����  oo/       Meeting     �5Z�U  P6Z�U  �-ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �2Z�U  ����  $p/      Workout     p;[�U  �;[�U  �<[This_stuffs_This_stuffs_ �U  p?[�U  �?[�U  p@[�U  �@[�U  ������  Nq/       Workout     &Z�U  �&Z�U  �'ZThis_stuffs_This_stuffs_ �U  P*Z�U  +Z�U  �+Z�U  �,Z�U  \�G���  ��/      Birthday    0�Z�U  �Z�U  ��ZThis_stuffs_This_stuffs_ �U  0�Z�U  �Z�U  p�Z�U  0�Z�U  �I����  H�/      Workout �U  p�Z�U  0�Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  ������  +�/       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             Խi���  ��/      Meeting �U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  yw���  J�/       Meeting     �WZ�U  @XZ�U   YZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `^Z�U  �x���  !/       Some_stuffs �Z�U  �Z�U  PZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Z�U  �����  4/      Meeting     5Y�U  �5Y�U  P8YSome_stuffs_Some_stuffs_ �U  @?Y�U  AY�U  EY�U  �EY�U  +V���  �/       Some_stuffs  �]�U  ��]�U   �]Some_stuffs_Some_stuffs_ �U  @�]�U  ��]�U  @�]�U  ��]�U  �����  �/       Workout     @�]�U  ��]�U  @�]This_stuffs_This_stuffs_ �U  @�]�U   �]�U  ��]�U  @�]�U  ����  _0/       Birthday    �[�U  P[�U  [justforfun_justforfun_ [�U  �[�U  �[�U  [�U  �[�U  \����  �0/      Appointment   Z�U  � Z�U  �!ZThis_stuffs_This_stuffs_ �U  �$Z�U  p-Z�U  &Z�U  �&Z�U  �q����  �0/       Birthday    PZ\�U  [\�U  �[\This_stuffs_This_stuffs_ �U  P^\�U  �^\�U  @�\�U  ��\�U  �7���  Z/       Workout �U  `]�U   ]�U  �]This_stuffs_This_stuffs_ �U  �]�U  @]�U    ]�U  � ]�U  �1����  ��/       Birthday nt ��]�U  p�]�U  ��]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��]�U  ������  �/      Appointment ��Z�U  ��Z�U  @�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `�Z�U  J.i���  =�/       Workout     �<Z�U  P=Z�U  >ZSome_stuffs_Some_stuffs_ �U  PAZ�U  �AZ�U  �BZ�U  PCZ�U  �9k���  è/       Birthday nt `Z�U   Z�U  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @Z�U  ��y���  z�/      Workout     ��Z�U  `�Z�U   �ZSome_stuffs_Some_stuffs_ �U  `�Z�U   �Z�U  ��Z�U  ��Z�U  :����  �/       Appointment  B^�U  �B^�U   C^justforfun_justforfun_ ^�U  `E^�U  F^�U  �F^�U  G^�U  �	���  /�/      Some_stuffs 0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  1����  ^�/       Some_stuffs �7\�U  P8\�U  �8\justforfun_justforfun_ \�U  �;\�U  P<\�U  �<\�U  �=\�U  x$����  ��/       Meeting     �0Z�U  p1Z�U  02ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �7Z�U  zq����  �/       Meeting     Pu[�U  �u[�U  Pv[This_stuffs_This_stuffs_ �U  �x[�U  �y[�U  ��[�U  p�[�U  �Ч���  ��/       Some_stuffs �+Z�U  �,Z�U  �5Zjustforfun_justforfun_ Z�U  0/Z�U  �/Z�U  �0Z�U  p1Z�U  �.����  ��/      Meeting ffs �\�U  ��\�U  �\justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  � ]�U  ��+���  �/      Meeting      �Y�U  ��Y�U  ��YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Z�U  ��,���  �/       Birthday    @p[�U   q[�U  �q[This_stuffs_This_stuffs_ �U  t[�U  �t[�U  Pu[�U  �u[�U  ��5���  $/       Birthday                       justforfun_justforfun_                                       3"6���  >/       Birthday    �[�U  `[�U   [Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �[�U  �%����  pF/       Birthday                       justforfun_justforfun_                                       ݣ����  [H/      Birthday     �\�U  ��\�U  ��\Some_stuffs_Some_stuffs_ �U  `�\�U   �\�U  ��\�U  `�\�U  I�Z���  i/       Appointment  �\�U  ��\�U  ��\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0�\�U  ��j���  4m/      Workout      �Y�U  ��Y�U  ��YSome_stuffs_Some_stuffs_ �U  P�Y�U  �Y�U  ��Y�U  ��Y�U  H�����  ]�/       Some_stuffs                    Some_stuffs_Some_stuffs_                                     �����  c�/      Some_stuffs `�\�U  ��\�U  ��\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��\�U  L����  A�/      Some_stuffs ��Y�U  ��Y�U  �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `�Y�U  Qp$���  R�/       Appointment �Z�U  �Z�U  `ZSome_stuffs_Some_stuffs_ �U  �Z�U  @Z�U    Z�U  � Z�U  H55���  ��/       Workout �U  xY�U  �xY�U  �|Yjustforfun_justforfun_ Y�U  ��Y�U  ��Y�U  p�Y�U  0�Y�U  &:���  ��/      Some_stuffs ��[�U  �[�U  ��[justforfun_justforfun_ \�U    \�U  � \�U  `\�U  �\�U  )"����  i/       Some_stuffs �x[�U  �y[�U  ��[Some_stuffs_Some_stuffs_ �U  �|[�U  p}[�U  0~[�U  �~[�U  d�����  @/      Birthday    p�Y�U  0�Y�U  0�Yjustforfun_justforfun_ Y�U   �Y�U  ��Y�U  ��Y�U  p�Y�U  ������  �/       Workout     �]�U  0]�U  �]This_stuffs_This_stuffs_ �U  0]�U  �]�U  0]�U  �]�U  �;s��  �#/       Meeting  U  �=]�U   >]�U  �>]justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  C]�U  �w��  !�#/       Appointment �]Z�U  `^Z�U   _ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `dZ�U  H~��  յ#/       Meeting     ��Y�U  ��Y�U  �Yjustforfun_justforfun_ Y�U  `�Y�U   �Y�U  ��Y�U  `�Y�U  �|��  $�#/       Meeting     �T]�U  �U]�U  V]justforfun_justforfun_ ]�U  �X]�U  �Y]�U  @Z]�U  �Z]�U  �{���  ��#/       Appointment �rZ�U  psZ�U  0tZSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  �xZ�U  <����  W�#/      Birthday U  �\�U  p\�U  0\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �\�U  �#��  �#/       Meeting �U  @�[�U  ��[�U  ��[justforfun_justforfun_ _This_stuffs_This_stuffs_ �U   �[�U  �Z*��  ��#/       Birthday nt 0�[�U  ��[�U  0�[This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  p�[�U  ̓-��  ��#/      Appointment �!Z�U  @"Z�U   #ZSome_stuffs_Some_stuffs_ �U  &Z�U  �&Z�U  �'Z�U  P(Z�U  |����  �$/      Workout     К]�U  P�]�U  Л]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��]�U  \�;��  �'$/      Some_stuffs @SZ�U   TZ�U  �TZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �YZ�U  ��@��  #)$/       Some_stuffs `�Z�U  �Z�U  `�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �Z�U  ��L��  C,$/       Meeting �U  Ш]�U  ��]�U   �]justforfun_justforfun_ ]�U  0�]�U  ��]�U  0�]�U  ��]�U  qPR��  �-$/       Birthday    p}Z�U  �}Z�U  �rZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  pwZ�U  �eU��  p.$/       Workout     @�\�U  ��\�U  �`\Some_stuffs_Some_stuffs_ �U  pc\�U  �c\�U  pd\�U  �d\�U  4�W��  �.$/       Birthday    P�[�U  ж[�U  P�[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  л[�U  �}���  �W$/      Some_stuffs �\]�U   ]]�U  �]]justforfun_justforfun_ ]�U  �_]�U  ``]�U  a]�U  �a]�U  ��x��  y$/       Birthday    ��X�U  ��X�U  0�Xjustforfun_justforfun_ X�U   �X�U  ��X�U  ��X�U  @�X�U  �b���  $/      Meeting     0�Z�U  ��Z�U  p�Zjustforfun_justforfun_ Z�U  ��Z�U  ��Z�U  0�Z�U  � [�U  �
��  �$/      Some_stuffs @�[�U  ��[�U  @�[This_stuffs_This_stuffs_ �U  ��[�U  @�[�U   �[�U  ��[�U  Ø��  ��$/       Some_stuffs @q]�U  �q]�U  @r]Some_stuffs_Some_stuffs_ �U  @t]�U  �t]�U  @u]�U   v]�U  !� ��  �$/       Meeting     �\�U  0\�U  �\justforfun_justforfun_ \�U  0\�U  �\�U  0\�U  �\�U  �,!��  $�$/       Appointment ��[�U  p�[�U  �[This_stuffs_This_stuffs_ �U  P�[�U  �[�U  ��[�U  �[�U  ����  9�$/       Some_stuffs                    This_stuffs_This_stuffs_                                     ����  ��$/       Appointment ��Y�U  ��Y�U  P�YThis_stuffs_This_stuffs_ �U  `�Y�U   �Y�U   �Y�U  ��Y�U  R�9 ��  ��$/       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             YBC ��  g�$/       Meeting     �QZ�U  �RZ�U  �HZThis_stuffs_This_stuffs_ �U  �KZ�U  pLZ�U  0MZ�U  �MZ�U  �bJ ��  :�$/      Some_stuffs �[�U  ��[�U  �[justforfun_justforfun_ [�U  ��[�U  �[�U  ��[�U  ��[�U  ��� ��  9%/       Meeting     �~]�U  @]�U   �]This_stuffs_This_stuffs_ �U  0�]�U  ��]�U   �]�U  ��]�U  ��� ��  :%/      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �T� ��  �%/       Appointment P�^�U  г^�U  ��^Some_stuffs_Some_stuffs_ �U  ж^�U  P�^�U  з^�U  ��^�U  q6h!��  f9%/       Workout     ��X�U  @�X�U   YSome_stuffs_Some_stuffs_ �U  PY�U  Y�U   	Y�U  �	Y�U  �u!��  �<%/      Birthday    ��[�U  `�[�U  �\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �\�U  P�x!��  �=%/       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             r��!��  A%/       Some_stuffs �Z�U  ��Z�U  @�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Z�U  ��"��  !h%/       Appointment  �]�U  ��]�U   �]This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  �]�U  d
�"��  @�%/      Appointment �\Z�U   ]Z�U  @SZThis_stuffs_This_stuffs_ �U  @VZ�U   WZ�U  �WZ�U  @XZ�U  ���"��  Í%/       Meeting     �Z�U  ��Z�U  0�Zjustforfun_justforfun_ Z�U  �Z�U  ��Z�U  @�Z�U  ��Z�U  �=#��  ��%/      Appointment �%Y�U  �&Y�U  )YSome_stuffs_Some_stuffs_ �U  �1Y�U  �2Y�U  5Y�U  �5Y�U  �z�#��  <�%/      Meeting �U   6_�U  �6_�U   7_justforfun_justforfun_ _�U   9_�U  �9_�U   :_�U  �:_�U  �8�#��  y�%/       Some_stuffs p?[�U  �?[�U  p@[justforfun_justforfun_ [�U  �B[�U  pC[�U  0D[�U  �D[�U  �c$��  ��%/       Some_stuffs ��[�U  @�[�U  ��[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��[�U  S�k$��  ��%/       Birthday     �]�U  ��]�U   �]Some_stuffs_Some_stuffs_ �U  ��]�U  `�]�U  ��]�U  `�]�U  ��q$��  � &/       Workout     Y\�U  �Y\�U  PZ\Some_stuffs_Some_stuffs_ �U   ]\�U  �]\�U  P^\�U  �^\�U  ��$��  �&/      Workout     P�[�U  �[�U  й[This_stuffs_This_stuffs_ �U  P�[�U  �[�U  н[�U  ��[�U  `<
%��  |'&/       Workout     ��Z�U  0�Z�U  �Zjustforfun_justforfun_ Z�U  ��Z�U  0�Z�U  �Z�U  ��Z�U  ���%��  Q&/      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �?&��  �v&/      Some_stuffs �zZ�U  �{Z�U  p|ZThis_stuffs_This_stuffs_ �U  �Z�U  ��Z�U  p�Z�U  0�Z�U  ��&��  ��&/       Appointment �$\�U  P%\�U  &\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  +\�U  �f�&��  �&/       Meeting     ��[�U   �[�U  ��[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @�[�U  <�`'��  ��&/      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             y2|'��  ��&/       Birthday    ��[�U  P�[�U  �[This_stuffs_This_stuffs_ �U  г[�U  ��[�U  �[�U  е[�U  $	�'��  ��&/      Birthday     \Z�U  pgZ�U  �]Zjustforfun_justforfun_ Z�U  �`Z�U  `aZ�U   bZ�U  �bZ�U  �9�(��  q'/      Appointment �Z�U  pZ�U  0	ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @Z�U  XG�(��  �'/       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ��(��  �'/       Some_stuffs �Y�U  `Y�U  �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �&Y�U  ��1)��  �7'/      Workout     P�Y�U  �Y�U  ��YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  4,�)��  �^'/      Meeting      ]\�U  �]\�U  P^\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �b\�U  P�a*��  ��'/       Some_stuffs ��X�U  @�X�U   YThis_stuffs_This_stuffs_ �U  PY�U  Y�U   	Y�U  �	Y�U  tci*��  ��'/       Workout �U  �_�U  P _�U  � _Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �$_�U  [�i*��  ��'/       Workout     p�Z�U  ��Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�Z�U  2�o*��  �'/       Meeting ent �w[�U  Px[�U  �x[This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  p}[�U  M�r*��  �'/      Workout �U  \�U  �\�U  @ \This_stuffs_This_stuffs_ �U  p"\�U  �"\�U  �#\�U  P$\�U  �zx*��  c�'/       Some_stuffs _�U  �_�U  @_Some_stuffs_Some_stuffs_ �U  p_�U   _�U  �_�U   _�U  ���*��  )�'/      Birthday      Z�U  � Z�U  �!ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �&Z�U  @^�*��  h�'/       Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             4R�+��  B�'/      Appointment 0�Z�U  �Z�U  p�ZSome_stuffs_Some_stuffs_ �U  �Z�U  ��Z�U  0�Z�U  �Z�U  i��+��  ��'/       Meeting ent ��\�U   �\�U  ��\This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  0�\�U  Y@W��  '�2/       Meeting ffs P4\�U  �4\�U  P5\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �9\�U  ��+W��  ��2/      Meeting     �Z�U  @Z�U  PZjustforfun_justforfun_ Z�U  PZ�U  �Z�U  �Z�U  PZ�U  	p�W��  �3/       Birthday    ��[�U  0�[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0�[�U  ظ�W��  w!3/       Some_stuffs ��Z�U   �Z�U   �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `�Z�U  {3�W��  ["3/       Birthday    �\�U  ��\�U  �\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��\�U  B�W��  �$3/      Meeting     �%Y�U  �&Y�U  )YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �5Y�U  ��CX��  �D3/      Birthday U  0MZ�U  �MZ�U  pNZThis_stuffs_This_stuffs_ �U  �\Z�U   ]Z�U  @SZ�U   TZ�U  �KX��  �F3/       Birthday U   eZ�U  �eZ�U  �fZThis_stuffs_This_stuffs_ �U  0iZ�U  �iZ�U  �jZ�U  pkZ�U  ��UX��  6I3/       Workout     �^�U  �^�U  `^Some_stuffs_Some_stuffs_ �U  �^�U  `^�U  �^�U  �^�U  8}�X��  �m3/       Some_stuffs @�\�U  ��\�U  @�\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��\�U  !b|Y��  ��3/       Meeting     �Z�U  �%Z�U  �ZThis_stuffs_This_stuffs_ �U  �!Z�U  @"Z�U   #Z�U  �#Z�U  ���Y��  G�3/      Appointment ��Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �Z�U  �q
Z��  �3/      Meeting     ��[�U   �[�U  ��[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @�[�U  �Z��  L�3/       Appointment �Y�U  `Y�U  �YSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  `#Y�U  �,Z��  v�3/       Workout     @VZ�U   WZ�U  �WZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  pgZ�U  ��Z��  ��3/       Workout     �e[�U   f[�U  �f[justforfun_justforfun_ [�U  @i[�U  �i[�U  @j[�U  �j[�U  S�'Z��  r�3/       Meeting     �PY�U  @QY�U  0TYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0bY�U  .!�Z��  ��3/      Workout     �gZ�U  phZ�U  0iZjustforfun_justforfun_ Z�U  0lZ�U  �lZ�U  pmZ�U  0nZ�U  ��Z��  J�3/       Meeting                        justforfun_justforfun_ _                                     �l�Z��  v�3/       Some_stuffs �[�U  p�[�U  0�[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �[�U  �K�Z��  ��3/       Meeting     `[�U   [�U  �[Some_stuffs_Some_stuffs_ �U  `	[�U   
[�U  �
[�U   [�U  �lB[��  �4/       Meeting     EY�U  �EY�U  �HYThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   VY�U  �DH[��  O
4/       Some_stuffs ��]�U  `�]�U  ��]justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  ��]�U  �'T[��  Z4/      Meeting     ��Z�U  ��Z�U  0�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `�Z�U  l��[��  U34/      Some_stuffs ��\�U  @�\�U  ��\justforfun_justforfun_ \�U  ��\�U  @�\�U  ��\�U  ��\�U  ��k\��  �T4/      Some_stuffs  �Y�U  �Y�U  0�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Y�U  ��n\��  �U4/       Meeting     �G\�U  PH\�U  �H\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �L\�U  [vs\��  �V4/       Some_stuffs �$]�U  p%]�U  �%]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �)]�U  �|}\��  xY4/       Workout     ��\�U  @�\�U  ��\This_stuffs_This_stuffs_ �U  p�\�U  �\�U  ��\�U   �\�U  �]��  �{4/      Meeting     �x\�U  @y\�U  �y\Some_stuffs_Some_stuffs_ �U   |\�U  �|\�U  @}\�U  �}\�U  8
]��  }4/       Meeting     �eY�U  `fY�U  �iYjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  �xY�U  �!]��  Y�4/       Appointment  �]�U  ��]�U   �]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �]�U  �¾]��  ��4/       Appointment  �Y�U  �Y�U  0�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Y�U  ��4^��  ��4/       Workout     �Z�U  �Z�U  `Zjustforfun_justforfun_ Z�U  �Z�U  @Z�U    Z�U  � Z�U  %�B^��  x�4/      Birthday    )Z�U  �)Z�U  P*ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �.Z�U  ���^��  ��4/      Some_stuffs                    Some_stuffs_Some_stuffs_                                     	��^��  ��4/       Workout      [�U  �[�U  `[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   
[�U  ��i_��  5/       Workout     �[�U  ��[�U  �[Some_stuffs_Some_stuffs_ �U  ��[�U  ��[�U  �[�U  ��[�U  $|�_��  �5/      Birthday    ��X�U  @�X�U   YThis_stuffs_This_stuffs_ �U  PY�U  Y�U   	Y�U  �	Y�U  J�_��  =?5/       Meeting ent  �Y�U  ��Y�U  ��YSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  �Z�U  �*`��  �A5/      Meeting �U  ��Y�U  ��Y�U  p�Yjustforfun_justforfun_ _ �U  p�Y�U  0�Y�U  ��Y�U  �Y�U  �``��  yE5/       Appointment `[�U  �[�U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P[�U  <)�`��  wg5/      Some_stuffs                    justforfun_justforfun_                                       �˱`��  m5/       Meeting ffs �1Y�U  �2Y�U  5YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  AY�U  ĽBa��  �5/      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             	rJa��  �5/       Some_stuffs `�Y�U   �Y�U   �Yjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ��Y�U  ��La��  ��5/       Appointment `�^�U  ��^�U  `�^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �^�U  �V�a��  �5/       Workout     @(]�U  �(]�U  p)]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   -]�U  ���a��  Q�5/      Appointment �vZ�U  pwZ�U  0xZSome_stuffs_Some_stuffs_ �U  �zZ�U  �{Z�U  p|Z�U  �|Z�U  3�a��  �5/       Birthday nt ��]�U  ��]�U   �]justforfun_justforfun_ _ his_stuffs_This_stuffs_ �U  ��]�U  {�a��  ��5/       Workout      �Y�U  �Y�U  0�YThis_stuffs_This_stuffs_ �U  ��Y�U  ��Y�U  P�Y�U  �Y�U  ��gb��  �5/      Workout �U  �jZ�U  pkZ�U  0lZjustforfun_justforfun_ Z�U  �nZ�U  �oZ�U  ppZ�U  0qZ�U  �c��  �6/       Meeting     �Z�U  �Z�U  PZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Z�U  �lc��  S	6/      Appointment �Z�U  @Z�U  PZSome_stuffs_Some_stuffs_ �U  PZ�U  �Z�U  �Z�U  PZ�U  ��c��  �-6/       Meeting ffs ��]�U  P�]�U  Ч]This_stuffs_This_stuffs_ �U   �]�U  ��]�U  0�]�U  ��]�U  Y�c��  �06/       Some_stuffs 0K[�U  �K[�U  c[Some_stuffs_Some_stuffs_ �U  pO[�U  �O[�U  pP[�U  0Q[�U  (�c��  �06/      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             e\.d��  �Q6/      Meeting     @SZ�U   TZ�U  �TZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �YZ�U  ��;d��  �T6/       Birthday    �TZ�U  �UZ�U  @VZSome_stuffs_Some_stuffs_ �U   YZ�U  �YZ�U  �ZZ�U  @[Z�U  ��Ld��  KY6/       Appointment 0�Z�U  ��Z�U  `�Zjustforfun_justforfun_ Z�U  @�Z�U   �Z�U  ��Z�U  ��Z�U  ��d��  Zy6/       Workout      �Y�U  ��Y�U  ��YThis_stuffs_This_stuffs_ �U  �Z�U  `Z�U   Z�U  �Z�U  0��d��  �z6/       Birthday                       This_stuffs_This_stuffs_                                     ���d��  $|6/       Appointment ��Z�U  0�Z�U  ��Zjustforfun_justforfun_ [�U  `�Z�U  ��Z�U  `�Z�U   �Z�U  %/�d��  �|6/      Birthday    p�Z�U  0�Z�U  ��ZThis_stuffs_This_stuffs_ �U  ��Z�U  ��Z�U  p�Z�U  ��Z�U  �]e��  .�6/      Some_stuffs L]�U  �L]�U  M]Some_stuffs_Some_stuffs_ �U  PO]�U  �O]�U  PP]�U  �P]�U  9^e��  J�6/       Birthday     �Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�Z�U  yWde��  ۠6/       Birthday    �A[�U  0B[�U  �B[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �G[�U  af��  ��6/       Workout     p�[�U  �[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��[�U  P>	f��  �6/       Appointment @�\�U  ��\�U  p�\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  Н\�U  ��f��  ��6/       Meeting     �C]�U  D]�U  �D]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0H]�U  ��f��  9�6/       Birthday    0�[�U  ��[�U  p�[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��[�U  |�Ag��  7/      Meeting     �[�U  е[�U  P�[This_stuffs_This_stuffs_ �U  P�[�U  �[�U  й[�U  ��[�U  �]h��  �c7/      Some_stuffs ��X�U  ��X�U  0�XThis_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  @�X�U  �'eh��  �e7/       Some_stuffs PO]�U  �O]�U  PP]Some_stuffs_Some_stuffs_ �U  �R]�U  pS]�U  �S]�U  pT]�U  :xqh��  �h7/       Birthday    �^�U  ��^�U  �^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��^�U  ��h��  <�7/      Meeting     P[�U  [�U  �[justforfun_justforfun_ [�U  �[�U  P[�U  �[�U  �[�U  ��i��  �7/       Appointment                    justforfun_justforfun_                                        l����  �;B/       Birthday    0]�U  �]�U  0]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0]�U  vA���  �^B/       Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �I���  �`B/      Some_stuffs �[�U  `[�U   [Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �[�U  �CL���  YaB/       Appointment @�[�U  ��[�U  @�[This_stuffs_This_stuffs_ �U  ��[�U  ��[�U   �[�U  ��[�U  �+ܓ��  0�B/      Birthday U  0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  �����  .�B/       Some_stuffs `�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �Z�U  6�p���  B�B/      Some_stuffs 0e_�U  �e_�U  0f_Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  �i_�U  q�p���  F�B/       Appointment �]�U  ��]�U  P�]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��]�U  ��x���  6�B/       Some_stuffs ��Y�U  ��Y�U  p�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  k���  ��B/      Appointment 1]�U  �1]�U  @2]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �5]�U  �w���  /�B/       Appointment ��Y�U  ��Y�U  �Yjustforfun_justforfun_ Y�U  `�Y�U   �Y�U  ��Y�U  `�Y�U  f����  `�B/      Workout �U  9^�U  �9^�U  p:^This_stuffs_This_stuffs_ �U  �<^�U  P=^�U  �=^�U  P>^�U  �\����  ��B/       Meeting     �9]�U  �:]�U   ;]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `?]�U  �����  C C/       Appointment �Z�U  ��Z�U   �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Z�U  2Q;���  �!C/       Some_stuffs 0�[�U  ��[�U  ��[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �[�U  �<���  
"C/       Appointment p�Z�U  0�Z�U  ��Zjustforfun_justforfun_ Z�U  0�Z�U  �Z�U  ��Z�U  0�Z�U  �xD���  �#C/       Some_stuffs p-[�U  �-[�U  �.[This_stuffs_This_stuffs_ �U  01[�U  �1[�U  �2[�U  03[�U  �K���  �%C/       Birthday U  �I]�U  �J]�U  K]Some_stuffs_Some_stuffs_ �U  M]�U  �M]�U  PN]�U  �N]�U  � X���  �(C/       Birthday      \�U  � \�U  `\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   \�U  �]���  l*C/       Appointment  �Y�U  ��Y�U  ��YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Z�U  ����  pLC/      Birthday nt ��Y�U  `�Y�U   �YThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ��Y�U  �o���  hpC/      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �;���  ,�C/       Workout     �jZ�U  pkZ�U  0lZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0qZ�U  �!���  .�C/      Birthday    `\�U   \�U  �\Some_stuffs_Some_stuffs_ �U   \�U  �\�U  `\�U   	\�U  ������  n�C/       Meeting     p�\�U  �\�U  p�\justforfun_justforfun_ \�U  ��\�U  p�\�U  �\�U  ��\�U  �ɲ���  F�C/      Meeting     �\�U  p\�U  0\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �\�U  Ȣ����  �C/       Workout     `�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_ �U   �Z�U  ��Z�U  `�Z�U  ��Z�U  B�=���  ��C/       Meeting ffs  �]�U  ��]�U   �]This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  `�]�U  �YN���  �C/       Some_stuffs  �Y�U  ��Y�U  ��YThis_stuffs_This_stuffs_ �U  ��Y�U  ��Y�U  �Y�U  ��Y�U  �hT���  ��C/      Appointment ��[�U  P�[�U  г[justforfun_justforfun_ [�U  P�[�U  ж[�U  P�[�U  з[�U  )hV���  )�C/       Birthday    �[�U  0�[�U  ��[This_stuffs_This_stuffs_ �U  p�[�U  0�[�U  ��[�U  0�[�U  �����  �D/       Meeting �U  ��Y�U  ��Y�U  p�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  u����  *D/      Workout     ��Y�U  ��Y�U  �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `�Y�U  ����  �D/       Workout ent P*Z�U  +Z�U  �+ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �/Z�U  �w���  D7D/      Meeting     5Y�U  �5Y�U  P8YThis_stuffs_This_stuffs_ �U  @?Y�U  AY�U  EY�U  �EY�U  ��}���  �8D/       Workout     ��Z�U  p�Z�U  0�ZSome_stuffs_Some_stuffs_ �U  ��Z�U  0�Z�U  ��Z�U  ��Z�U  :�����  �;D/       Meeting     p�Z�U  0�Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0�Z�U  �L#���  &cD/      Meeting     ��[�U  P�[�U  �[Some_stuffs_Some_stuffs_ �U  ��[�U  `�[�U   �[�U  ��[�U  1�����  ��D/       Some_stuffs ��Y�U  ��Y�U  p�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  <S����  ��D/      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �=����  A�D/       Workout �U  0\�U  �\�U  �\Some_stuffs_Some_stuffs_ �U  �\�U  p\�U  0\�U  �\�U  y7���  ۩D/       Birthday U  0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  �K���  ܮD/      Some_stuffs ��Y�U  ��Y�U  p�YThis_stuffs_This_stuffs_ �U  ��Y�U  @�Y�U   �Y�U  ��Y�U  $�ܜ��  8�D/      Some_stuffs �[�U  �[�U  [This_stuffs_This_stuffs_ �U  �[�U  �[�U  P[�U  [�U  �Ip���  ��D/       Workout     �V[�U  �W[�U  pX[Some_stuffs_Some_stuffs_ �U  0[[�U  �[[�U  0\[�U  �\[�U  eZy���  @�D/      Meeting     ��Y�U  ��Y�U  �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `�Y�U  XȀ���  '�D/       Meeting     ��Y�U  ��Y�U   �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  `���  �#E/       Meeting     ��Z�U  ��Z�U  @�ZThis_stuffs_This_stuffs_ �U   �Z�U  ��Z�U  ��Z�U   �Z�U  򳜞��  �FE/       Meeting     �+Z�U  �,Z�U  �5Zjustforfun_justforfun_ Z�U  0/Z�U  �/Z�U  �0Z�U  p1Z�U  ������  �GE/      Appointment ��Y�U  `�Y�U   �Yjustforfun_justforfun_ Y�U  p�Y�U  0�Y�U  ��Y�U  ��Y�U  �ӥ���  ,IE/       Meeting     �Y�U  @ Y�U  �"YThis_stuffs_This_stuffs_ �U  )Y�U  �)Y�U  p-Y�U  0.Y�U  �ǩ���  /JE/       Meeting �U  ��Z�U  p�Z�U  0�Zjustforfun_justforfun_ Z�U  ��Z�U  0�Z�U  �Z�U  ��Z�U  �SI���  sE/      Some_stuffs ��X�U  @�X�U   YThis_stuffs_This_stuffs_ �U  PY�U  Y�U   	Y�U  �	Y�U  ��K���  �sE/       Some_stuffs p@[�U  �@[�U  �A[justforfun_justforfun_ [�U  0D[�U  �D[�U  �E[�U  0F[�U  �#O���  �tE/       Workout                        This_stuffs_This_stuffs_                                     �ҟ��  *�E/       Appointment �\�U  p\�U  0\This_stuffs_This_stuffs_ �U  �\�U  p\�U  �\�U  p\�U  0�؟��  ��E/       Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �Oޟ��  +�E/       Some_stuffs �^]�U  `_]�U  �_]Some_stuffs_Some_stuffs_ �U  0b]�U  �b]�U  pc]�U  �c]�U  �3���  0�E/      Birthday    ��^�U   �^�U  ��^Some_stuffs_Some_stuffs_ �U  `�^�U  �^�U  `�^�U  �^�U  b�^���  ��E/       Workout     `4]�U  �4]�U  `5]justforfun_justforfun_ ]�U  �7]�U   8]�U  �8]�U  `9]�U  \Wl���  ��E/       Birthday    ��X�U  ��X�U  0�XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @�X�U  Q�p���  ��E/       Meeting     �>]�U  `?]�U  �?]This_stuffs_This_stuffs_ �U  `B]�U  C]�U  �C]�U  D]�U  �~���  D�E/      Workout     ��X�U  @�X�U   YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �	Y�U  c����  |�E/       Meeting     ��Y�U  ��Y�U  p�YThis_stuffs_This_stuffs_ �U  ��Y�U  @�Y�U   �Y�U  ��Y�U  rd����  &�E/       Some_stuffs ��Y�U  @�Y�U  ��YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  � Z�U  v	���  ��E/       Some_stuffs ��Y�U  ��Y�U  p�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Y�U  �����  ��E/       Some_stuffs                    justforfun_justforfun_                                       ����  ��E/      Some_stuffs �Z�U  @Z�U  PZSome_stuffs_Some_stuffs_ �U  PZ�U  �Z�U  �Z�U  PZ�U  �#0���  01F/       Some_stuffs ��[�U   �[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @�[�U  Ξ1���  �1F/      Workout ffs ��]�U   �]�U  ��]This_stuffs_This_stuffs_ �U   �]�U  ��]�U   �]�U  ��]�U  � D���  N6F/       Birthday    �[�U  �$[�U  �[justforfun_justforfun_ [�U  P[�U  [�U  �[�U  �[�U  o����  �UF/       Meeting     �[�U  0�[�U  ��[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0�[�U  T�Ţ��  rWF/       Workout     �m\�U   n\�U  �n\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @s\�U  "�ˢ��  YF/       Meeting     0�[�U  ��[�U  0�[This_stuffs_This_stuffs_ �U  ��[�U  p�[�U  �[�U  ��[�U  =�֢��  �[F/      Some_stuffs 0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  �ߢ��  ^F/       Meeting     ��Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_ �U  `�Z�U   �Z�U  ��Z�U  `�Z�U  1^���  ~~F/       Some_stuffs PQ]�U  ��]�U  �R]justforfun_justforfun_ ]�U  �T]�U  �U]�U  V]�U  �V]�U  0�z���  ޅF/       Some_stuffs p�Y�U  0�Y�U  0�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p�Y�U  ������  ץF/       Workout     оZ�U  P�Z�U  0�Zjustforfun_justforfun_ Z�U  0�Z�U  ��Z�U  0�Z�U  �Z�U  �>����  ��F/       Appointment �Z�U  ��Z�U   �ZSome_stuffs_Some_stuffs_ �U  оZ�U  P�Z�U  0�Z�U  �Z�U  46���  ¨F/      Workout ent                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             S���  �F/       Meeting     ��[�U  ��[�U  �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��[�U  �+K���  �{Q/      Meeting     0�Z�U  ��Z�U  p�Zjustforfun_justforfun_ Z�U  ��Z�U  ��Z�U  0�Z�U  � [�U  ������  Y�Q/       Some_stuffs �[�U  ��[�U  ��[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��[�U  \ku���  �Q/      Birthday U  0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��X�U  B����  ��Q/       Appointment 0)[�U  �)[�U  �*[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p/[�U  )	����  ��Q/       Birthday U  0~[�U  �~[�U  �[Some_stuffs_Some_stuffs_ �U  0�[�U  ��[�U  p�[�U  0�[�U  �<���  ~�Q/      Meeting                        justforfun_justforfun_                                       k���  ��Q/       Workout     p{[�U  0|[�U  �|[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�[�U  �$���  ��Q/       Birthday fs 0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  (�*���  i�Q/       Birthday nt P*\�U  +\�U  �+\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P0\�U  ������  DR/       Appointment                    Some_stuffs_Some_stuffs_                                     %����  xR/      Appointment p�Y�U  0�Y�U  0�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p�Y�U  �����  �hR/      Birthday    EY�U  �EY�U  �HYThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   VY�U  ������  lR/       Meeting �U  0~[�U  �~[�U  �[This_stuffs_This_stuffs_ �U  0�[�U  ��[�U  p�[�U  0�[�U  �x���  Q�R/      Appointment ��Z�U  ��Z�U  0�ZThis_stuffs_This_stuffs_ �U  `�Z�U   �Z�U  ��Z�U  `�Z�U  ����  ��R/      Some_stuffs                    justforfun_justforfun_                                       de����   �R/      Appointment 0TY�U   VY�U  @YYThis_stuffs_This_stuffs_ �U  paY�U  0bY�U  �eY�U  `fY�U  ��<���  .S/       Some_stuffs �rZ�U  psZ�U  0tZjustforfun_justforfun_ Z�U  �vZ�U  pwZ�U  0xZ�U  �xZ�U  ��<���  ;S/      Meeting �U  ��Z�U  ��Z�U  0�ZSome_stuffs_Some_stuffs_ �U  `�Z�U   �Z�U  ��Z�U  `�Z�U  TS���  �S/       Meeting      
^�U  �
^�U   ^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �^�U  H�����  )S/       Meeting     �Z�U  pZ�U  0	Zjustforfun_justforfun_ Z�U  �Z�U  �Z�U  �Z�U  @Z�U  �U����  �.S/      Appointment p�\�U  ��\�U  ��\This_stuffs_This_stuffs_ �U  ��\�U  @�\�U   �\�U  ��\�U  �����  �/S/       Some_stuffs PM\�U  �M\�U  PN\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  PR\�U  ��u���  [QS/      Birthday      Z�U  � Z�U  �!Zjustforfun_justforfun_ Z�U  �$Z�U  p-Z�U  &Z�U  �&Z�U  2}���  @SS/       Appointment  �\�U  ��\�U   �\This_stuffs_This_stuffs_ �U  ��\�U   �\�U  ��\�U   �\�U  ",���  �vS/       Some_stuffs �[�U  �$[�U  �[justforfun_justforfun_ [�U  P[�U  [�U  �[�U  �[�U  !���  xS/       Birthday    ��X�U  @�X�U   YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �	Y�U  �l#���  �}S/       Meeting     @oY�U   pY�U  �sYThis_stuffs_This_stuffs_ �U  �|Y�U  P}Y�U   �Y�U  ��Y�U  tQ%���  J~S/      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ԡ���  *�S/       Workout     ��Y�U  ��Y�U   �Yjustforfun_justforfun_ Y�U  ��Y�U  ��Y�U   �Y�U  ��Y�U  �����  ��S/       Appointment 0�Z�U  ��Z�U  0�ZSome_stuffs_Some_stuffs_ �U  ��Z�U  0�Z�U  �Z�U  ��Z�U  $����  ��S/       Appointment ��[�U  P�[�U  �[justforfun_justforfun_ [�U  ��[�U  `�[�U  �\�U  P\�U  6C����  �S/      Appointment  YZ�U  �YZ�U  �ZZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �_Z�U  hk����  ��S/       Birthday U  0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��X�U  j�8���  ��S/       Birthday fs 0�^�U  ��^�U  ��^Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  ��^�U  6;���  n�S/      Meeting     puZ�U  0vZ�U  �vZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �{Z�U  ��T���  ��S/       Some_stuffs �BZ�U  PCZ�U  DZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �RZ�U  ������  ��S/       Some_stuffs ��Y�U  ��Y�U  �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @�Y�U  �����  ��S/      Some_stuffs ��\�U  `�\�U  ��\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @�\�U  �\|���  �T/       Birthday    p3Z�U  04Z�U  �4ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P:Z�U  �����  (?T/      Meeting      �[�U  ��[�U  ��[This_stuffs_This_stuffs_ �U  ��[�U  �[�U  ��[�U  ��[�U  �K����  �dT/       Birthday    �^�U  ��^�U  �^This_stuffs_This_stuffs_ �U  ��^�U   �^�U  ��^�U   �^�U  �eL���  p�T/       Appointment                    justforfun_justforfun_                                       x����  ۭT/       Appointment `_^�U  ��^�U  ``^justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  d^�U  ��l���  E�T/      Some_stuffs �~Z�U  0Z�U  �ZThis_stuffs_This_stuffs_ �U  ��Z�U  ��Z�U  p�Z�U  0�Z�U  �.q���  d�T/       Appointment @�\�U  ��\�U  @�\justforfun_justforfun_ _ �U  `�\�U   �\�U  ��\�U   �\�U  �\w���  ��T/       Meeting  fs 0�[�U  ��[�U  ��[This_stuffs_This_stuffs_ �U  0�[�U  ��[�U  ��[�U  0�[�U  ������  C#U/       Birthday    p�Y�U  0�Y�U  0�YThis_stuffs_This_stuffs_ �U   �Y�U  ��Y�U  ��Y�U  p�Y�U  ������  �'U/      Appointment ��Y�U  `�Y�U   �Yjustforfun_justforfun_ Y�U  p�Y�U  0�Y�U  ��Y�U  ��Y�U  �-���  %KU/      Meeting     �'[�U  p([�U  0)[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �-[�U  �3���  �LU/       Some_stuffs `�Y�U   �Y�U   �YThis_stuffs_This_stuffs_ �U  p�Y�U  0�Y�U  ��Y�U  ��Y�U  ������  �xU/       Workout     �QZ�U  �RZ�U  �HZSome_stuffs_Some_stuffs_ �U  �KZ�U  pLZ�U  0MZ�U  �MZ�U  H����  �xU/       Workout      �\�U  ��\�U  ��\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0�\�U  �c���  �U/       Some_stuffs ��[�U  P�[�U  �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �[�U  �]{���  ��U/      Birthday    �<Z�U  P=Z�U  >Zjustforfun_justforfun_ Z�U  PAZ�U  �AZ�U  �BZ�U  PCZ�U  �����  )�U/      Meeting     ��Z�U  0�Z�U  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  ]����  +�U/      Workout     ��Y�U  ��Y�U  �Yjustforfun_justforfun_ Y�U  `�Y�U   �Y�U  ��Y�U  `�Y�U  ������  0�U/       Some_stuffs 0�[�U  ��[�U  0�[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��[�U  �v<���  �V/      Appointment  �Y�U  ��Y�U  ��YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Z�U  )G���  IV/       Appointment ��Y�U  ��Y�U  p�YThis_stuffs_This_stuffs_ �U  ��Y�U  @�Y�U   �Y�U  ��Y�U  D��	��  l�`/      Appointment                    justforfun_justforfun_                                       M}
��  ��`/      Appointment P:\�U  ;\�U  �;\justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  @?\�U  �h~
��  ��`/       Birthday    0�[�U  �[�U  ��[justforfun_justforfun_ [�U  0�[�U  ��[�U  p�[�U  0�[�U  ���
��  ��`/       Some_stuffs ��^�U   �^�U  ��^This_stuffs_This_stuffs_ �U  �_�U  `_�U  _�U  �_�U  �,��  �a/      Birthday U  �BZ�U  PCZ�U  DZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �RZ�U  ��,��  �a/       Meeting     ��Y�U  ��Y�U  p�Yjustforfun_justforfun_ Y�U  ��Y�U  @�Y�U   �Y�U  ��Y�U  �����  /5a/       Appointment `�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_ �U  `�Z�U   �Z�U  ��Z�U  ��Z�U  ����  :5a/       Some_stuffs �[�U  �[�U  `[justforfun_justforfun_ [�U   [�U  �[�U  �[�U  �$[�U  3Y���  �6a/       Meeting     �eY�U  `fY�U  �iYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �xY�U  �����  �7a/       Meeting �U  ��Y�U  `�Y�U   �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  ����  �9a/       Birthday                       Some_stuffs_Some_stuffs_                                     9R��  �\a/       Meeting     ��Y�U  p�Y�U  ��Yjustforfun_justforfun_ Y�U  �Y�U  ��Y�U   �Y�U  �Y�U  ,�_��  -`a/      Some_stuffs �Z�U  @Z�U  PZSome_stuffs_Some_stuffs_ �U  PZ�U  �Z�U  �Z�U  PZ�U  HM���  ��a/       Workout     P�^�U  к^�U  P�^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �^�U  �s���  ��a/      Birthday fs �_�U  `_�U  �_Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  `_�U  ����  �a/      Workout     �w\�U   x\�U  �x\justforfun_justforfun_ \�U   {\�U  �{\�U   |\�U  �|\�U  m���  �a/      Meeting     �<Z�U  P=Z�U  >Zjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  PCZ�U  ��!��  Y�a/       Appointment  �Y�U  �Y�U  0�Yjustforfun_justforfun_ Y�U  ��Y�U  ��Y�U  P�Y�U  �Y�U  |z���  ��a/      Birthday    ��Z�U  ` [�U  `[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   [�U  I����  ��a/       Meeting     `\�U   \�U  �\justforfun_justforfun_ \�U   \�U  �\�U  `\�U   	\�U  �*B��  :b/       Birthday    �W\�U  PX\�U  Y\This_stuffs_This_stuffs_ �U  �[\�U  P\\�U   ]\�U  �]\�U  �L��  �b/       Birthday    �/^�U   0^�U  �0^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   5^�U  ,	T��  �!b/      Appointment ��X�U  ��X�U  0�XThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @�X�U  :W��  �"b/       Birthday    �cZ�U  `dZ�U   eZjustforfun_justforfun_ _ �U  �gZ�U  phZ�U  0iZ�U  �iZ�U  y!Y��  #b/       Appointment �B\�U  @C\�U   D\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  PH\�U  �r��  kb/       Appointment @�[�U   �[�U   �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �[�U  \u���  Krb/      Meeting ffs �w[�U  Px[�U  �x[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p}[�U  �w"��  /�b/       Workout ent ��\�U  0�\�U  ��\This_stuffs_This_stuffs_ �U  ��\�U  `�\�U  �\�U  ��\�U  `���  \�b/       Some_stuffs 0MZ�U  �MZ�U  pNZjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U   TZ�U  #[���  4�b/       Birthday    �_\�U  `\�U  �>\Some_stuffs_Some_stuffs_ �U  @A\�U   B\�U  �B\�U  @C\�U  Y����  '�b/       Some_stuffs ��Z�U  `�Z�U   �ZThis_stuffs_This_stuffs_ �U  ��Z�U  ��Z�U  0�Z�U  ��Z�U  D����  (�b/       Appointment ��]�U  p�]�U  ��]justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  ��]�U  np���  վb/      Some_stuffs �U[�U  0V[�U  �V[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �[[�U  :��  ��b/       Meeting     �^�U   ^�U  �^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �^�U  !�<��  t�b/       Workout     ��Z�U   �Z�U   �ZSome_stuffs_Some_stuffs_ �U  `�Z�U   �Z�U  ��Z�U  `�Z�U  ��<��  ��b/       Appointment �[\�U  P\\�U   ]\justforfun_justforfun_ _ �U  @�\�U  ��\�U  �`\�U  0a\�U  ��G��  M�b/       Workout     PZ�U  Z�U  �ZThis_stuffs_This_stuffs_ �U  �Z�U  PZ�U  Z�U  �Z�U  
'���  5c/       Appointment ��X�U  @�X�U   YThis_stuffs_This_stuffs_ �U  PY�U  Y�U   	Y�U  �	Y�U  ty���  Jc/      Workout �U  0TY�U   VY�U  @YYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `fY�U  �����  �	c/       Meeting ent p�]�U  ��]�U  p�]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�]�U  �����  �
c/       Appointment  �Y�U  ��Y�U  ��YSome_stuffs_Some_stuffs_ �U  P�Y�U  �Y�U  ��Y�U  ��Y�U  ��r��  �/c/       Workout                        This_stuffs_This_stuffs_                                     �nt��  =0c/      Birthday    �eY�U  `fY�U  �iYjustforfun_justforfun_ Y�U  �sY�U  `tY�U  xY�U  �xY�U  ����  95c/       Meeting      	Y�U  �	Y�U  �YThis_stuffs_This_stuffs_ �U  �Y�U  `Y�U  �Y�U  `Y�U  4���  �[c/      Appointment p3Z�U  04Z�U  �4Zjustforfun_justforfun_ _This_stuffs_This_stuffs_ �U  P:Z�U  �P���  �~c/       Appointment puZ�U  0vZ�U  �vZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �{Z�U  d�B��  ��c/      Meeting     �eY�U  `fY�U  �iYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �xY�U  BG��  ��c/       Meeting      	Y�U  �	Y�U  �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `Y�U  �����  �c/       Appointment �[�U  P[�U  [This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �[�U   ����  ��c/       Appointment                    justforfun_justforfun_                                       �����  ��c/       Workout     7Z�U  �7Z�U  P8ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P=Z�U  �d��  ��c/      Some_stuffs 0TY�U   VY�U  @YYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `fY�U  �.��  �d/      Birthday    @SZ�U   TZ�U  �TZThis_stuffs_This_stuffs_ �U  �WZ�U  @XZ�U   YZ�U  �YZ�U  ���  yd/       Workout     �]�U  0]�U  �]justforfun_justforfun_ ]�U  0]�U  �]�U  p]�U  0]�U  �z���  >Ed/      Workout �U  �%Y�U  �&Y�U  )YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �5Y�U  �F���  7Fd/       Birthday    ��Y�U  ��Y�U  P�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  ����  nFd/       Meeting     0\[�U  �\[�U  �][Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0b[�U  v.��  �ed/      Some_stuffs `^�U   ^�U  �^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �^�U  ��5��  �gd/       Appointment �%Y�U  �&Y�U  )YThis_stuffs_This_stuffs_ �U  �1Y�U  �2Y�U  5Y�U  �5Y�U  �>M��  �md/       Meeting ffs �<\�U  �=\�U  �_\This_stuffs_This_stuffs_ �U  �?\�U  �@\�U  @A\�U   B\�U  �����  ��d/      Birthday    �eY�U  `fY�U  �iYThis_stuffs_This_stuffs_ �U  �sY�U  `tY�U  xY�U  �xY�U  �+���  ,�d/       Workout     ��Y�U  ��Y�U  p�Yjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ��Y�U  �d��  C�d/       Meeting      �Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   [�U  �nw��  9�d/       Meeting     �3[�U  p4[�U  �4[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pM[�U  9���  ��d/       Meeting     �\�U  ��\�U  @�\This_stuffs_This_stuffs_ �U  ��\�U   �\�U  ��\�U  @�\�U  8���  ��d/       Appointment �|]�U   }]�U  �}]Some_stuffs_Some_stuffs_ �U   �]�U  ��]�U  0�]�U  ��]�U  �_���  �e/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ����  te/      Meeting ent L\�U  �L\�U  PM\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  PQ\�U  �,��  %*e/      Birthday    ��Y�U  @�Y�U  ��Yjustforfun_justforfun_ Y�U  ��Y�U  `�Y�U    Z�U  � Z�U  U�wE��  ��o/      Workout �U  @l\�U  �l\�U  �m\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   r\�U  B�zE��  ��o/       Meeting     �/^�U   0^�U  �0^This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U   5^�U   ��E��   p/       Some_stuffs 0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��X�U  �dF��  z%p/       Meeting     P�[�U  п[�U  ��[Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  ��[�U  @5#F��  �)p/       Birthday                       Some_stuffs_Some_stuffs_                                     ��(F��  A+p/       Some_stuffs 0�Z�U  �Z�U  ��Zjustforfun_justforfun_ _ �U  @�Z�U  ��Z�U  �Z�U  p�Z�U  �1F��  �-p/       Meeting     @i[�U  �i[�U  @j[This_stuffs_This_stuffs_ �U  �l[�U   m[�U  �m[�U  �n[�U  m2F��  �-p/      Appointment `�Y�U   �Y�U   �YThis_stuffs_This_stuffs_ �U  p�Y�U  0�Y�U  ��Y�U  ��Y�U  h��F��  QPp/       Some_stuffs ��X�U  @�X�U   YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �	Y�U  ~�F��  �Pp/      Some_stuffs �Y�U  @ Y�U  �"YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0.Y�U  � ]G��  %zp/      Appointment  eZ�U  �eZ�U  �fZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pkZ�U  �R�G��  >�p/      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             *e�G��  I�p/       Workout     p]�U  �]�U  p]justforfun_justforfun_ ]�U  �]�U  0]�U  �]�U  �]�U  ��G��  ˠp/       Workout     �Z�U  ��Z�U   �ZSome_stuffs_Some_stuffs_ �U  оZ�U  P�Z�U  0�Z�U  �Z�U  ��{H��  ��p/      Meeting     ��Y�U  ��Y�U  p�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  aI��  ��p/       Appointment оZ�U  P�Z�U  0�ZSome_stuffs_Some_stuffs_ �U  0�Z�U  ��Z�U  0�Z�U  �Z�U  �I��  T�p/      Some_stuffs ��Y�U  ��Y�U  p�YSome_stuffs_Some_stuffs_ �U  p�Y�U  0�Y�U  ��Y�U  �Y�U   �&I��  T�p/       Birthday    ��Y�U  @�Y�U  ��YSome_stuffs_Some_stuffs_ �U  ��Y�U  @�Y�U  ��Y�U  ��Y�U  �#.I��  0�p/       Birthday    ��\�U  `�\�U   �\This_stuffs_This_stuffs_ �U  ��\�U  `�\�U  ��\�U  `�\�U  r�I��  Dq/      Workout      YZ�U  �YZ�U  �ZZThis_stuffs_This_stuffs_ �U  �]Z�U  `^Z�U   _Z�U  �_Z�U  ���I��  �q/       Birthday    P[�U  [�U  �[justforfun_justforfun_ [�U   [�U  � [�U  P![�U  "[�U  `'�I��  \q/       Workout                        justforfun_justforfun_                                       �SJ��  L<q/       Meeting     �B\�U  @C\�U   D\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  PH\�U  ��SJ��  O<q/       Appointment �
[�U   [�U  �[justforfun_justforfun_ [�U  �[�U  `[�U   [�U  �[�U  !�SJ��  T<q/       Some_stuffs 0�Z�U  ��Z�U  ��ZThis_stuffs_This_stuffs_ �U  p�Z�U  0�Z�U  ��Z�U  p�Z�U  ��XJ��  �=q/      Some_stuffs ��X�U  @�X�U   YThis_stuffs_This_stuffs_ �U  PY�U  Y�U   	Y�U  �	Y�U  "`_J��  T?q/       Appointment ��\�U  P�\�U  ��\Some_stuffs_Some_stuffs_ �U  �\�U  ��\�U  ��\�U   �\�U  ���J��  +_q/       Appointment 0�[�U  ��[�U  ��[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0�[�U  ���J��  (`q/      Appointment ��\�U  `�\�U   �\Some_stuffs_Some_stuffs_ �U  `�\�U  ��\�U  ��\�U  p$]�U  x��J��  {aq/       Birthday U  &Z�U  �&Z�U  �'ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �,Z�U  ���K��  Z�q/       Some_stuffs �eY�U  `fY�U  �iYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �xY�U  ��K��  j�q/       Birthday U  `�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_ �U  `[�U   [�U  �[�U  `[�U  �x�K��  ��q/       Workout                        Some_stuffs_Some_stuffs_                                     `YL��  ��q/       Some_stuffs @oY�U   pY�U  �sYThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  QCL��  2�q/       Some_stuffs p�Z�U  0�Z�U  ��ZThis_stuffs_This_stuffs_ �U  ��Z�U  ��Z�U  p�Z�U  ��Z�U  .�!L��  ��q/      Meeting      eZ�U  �eZ�U  �fZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  pkZ�U  ���L��  ��q/      Appointment                    justforfun_justforfun_                                       (a�L��  ��q/       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             l�L��  ��q/       Some_stuffs ��X�U  ��X�U  0�XThis_stuffs_This_stuffs_ �U   �X�U  ��X�U  ��X�U  @�X�U  #[�L��  4�q/       Birthday    �[�U  е[�U  P�[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��[�U  ���L��  b�q/       Workout      �Y�U  �Y�U  0�YThis_stuffs_This_stuffs_ �U  ��Y�U  ��Y�U  P�Y�U  �Y�U  )SHM��  	�q/       Some_stuffs ��\�U  ��\�U  @�\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �\�U  <JM��  w�q/      Birthday nt �,\�U  P-\�U  .\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �2\�U  t��M��  
#r/      Some_stuffs p�Y�U  0�Y�U  0�Yjustforfun_justforfun_ Y�U   �Y�U  ��Y�U  ��Y�U  p�Y�U  2-�M��  #r/       Birthday U  �]�U   ]�U  �]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �!]�U  ���M��  �%r/       Appointment `�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_ �U  `�Z�U   �Z�U  �Z�U  `�Z�U  9jN��  3Hr/       Some_stuffs ��Y�U  ��Y�U  �YThis_stuffs_This_stuffs_ �U  `�Y�U   �Y�U  ��Y�U  `�Y�U  ��wN��  �Kr/      Workout     �nZ�U  �oZ�U  ppZjustforfun_justforfun_ Z�U  �rZ�U  psZ�U  0tZ�U  �tZ�U  �~O��  rr/       Meeting     p%[�U  0&[�U  �&[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p+[�U  ��O��  $sr/       Meeting     p|Z�U  �|Z�U  �~Zjustforfun_justforfun_ Z�U  p�Z�U  0�Z�U  ��Z�U  ��Z�U  �O��  ��r/       Some_stuffs @�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �Z�U  ql�O��  &�r/       Meeting �U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��X�U  ��O��  %�r/       Workout                        Some_stuffs_Some_stuffs_                                     �?�O��  ��r/      Workout     �;Y�U  `<Y�U  @?Yjustforfun_justforfun_ Y�U  �HY�U  �IY�U  �LY�U  `MY�U  y�2P��  �r/       Appointment P'\�U  (\�U  �(\Some_stuffs_Some_stuffs_ �U  �+\�U  P,\�U  �,\�U  P-\�U  �BP��  C�r/      Some_stuffs ��[�U   �[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @�[�U  e�P��  ��r/       Some_stuffs 0 ]�U  � ]�U  0]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p]�U  �?�P��  Z�r/      Some_stuffs ��Y�U  ��Y�U  �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `�Y�U  �Q��  �s/       Meeting      �Y�U  �Y�U  0�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Y�U  �^�Q��  s/       Appointment @k[�U  �k[�U  �l[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   q[�U  ��R��  �6s/       Some_stuffs p-[�U  �-[�U  �.[This_stuffs_This_stuffs_ �U  01[�U  �1[�U  �2[�U  03[�U  %�R��  87s/      Meeting �U   �\�U  ��\�U  ��\justforfun_justforfun_ \�U  ��\�U  0�\�U  ��\�U  0�\�U  �R��  d\s/      Some_stuffs p�Z�U  ��Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Z�U  �MS��  z�s/       Workout     �n\�U  @o\�U  �o\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �t\�U  k�S��  ��s/      Appointment p�\�U  �\�U  ��\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @�\�U  ��S��  l�s/       Meeting     ��\�U  ��\�U  0�\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�\�U  �$rT��  ~�s/      Appointment ��Y�U  ��Y�U   �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  �$	U��  &�s/      Appointment  [�U  �[�U  `	[justforfun_justforfun_ _ �U  �[�U  �[�U  `[�U  �[�U  H��U��  ]t/       Workout     @�Z�U  ��Z�U  ��ZSome_stuffs_Some_stuffs_ �U  ��Z�U   �Z�U   �Z�U  ��Z�U  t��U��  & t/       Birthday     �Y�U  �Y�U  0�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Y�U  ���U��  E!t/       Meeting     �\�U  p\�U  �\Some_stuffs_Some_stuffs_ �U  @ \�U  � \�U  @!\�U  �!\�U  ��U��  �$t/      Appointment ��[�U  ��[�U  @�[justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  ��[�U  !ܯU��  �$t/       Workout ffs ��\�U  `�\�U   �\This_stuffs_This_stuffs_ �U  ��\�U  �\�U  ��\�U  0�\�U  ��,V��  �Dt/      Some_stuffs ��Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U   �Z�U  9�CV��  �Jt/       Some_stuffs P*\�U  +\�U  �+\Some_stuffs_Some_stuffs_ �U  .\�U  �.\�U  �/\�U  P0\�U  ȕHV��  �Kt/       Meeting     �8\�U  �9\�U  P:\justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  `\�U  �KV��  �Lt/       Appointment ��]�U  �]�U  ��]This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ^�U  ��V��  Znt/      Workout     �_\�U  `\�U  �>\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @C\�U  ���V��  pt/       Appointment �Z�U  ��Z�U  p�ZThis_stuffs_This_stuffs_ �U  0�Z�U  ��Z�U  @�Z�U   �Z�U  ���V��  Yst/       Birthday    �HZ�U  �IZ�U  0JZSome_stuffs_Some_stuffs_ �U  0MZ�U  �MZ�U  pNZ�U  0OZ�U  ٮnW��  7�t/       Meeting     ��Y�U  ��Y�U  p�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  �>uW��  �t/       Some_stuffs 7Z�U  �7Z�U  P8ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P=Z�U  L!"���  !D/      Some_stuffs �"[�U  #[�U  �#[This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  p([�U  �)6���  BI/       Meeting      �Y�U  ��Y�U  ��YSome_stuffs_Some_stuffs_ �U  ��Y�U  ��Y�U  �Y�U  ��Y�U  b����  Dg/      Appointment ��Z�U  `�Z�U   �ZThis_stuffs_This_stuffs_ �U  ��Z�U  `�Z�U  ��Z�U  ` [�U  �C���  J�/       Some_stuffs �<Z�U  P=Z�U  >ZSome_stuffs_Some_stuffs_ �U  PAZ�U  �AZ�U  �BZ�U  PCZ�U  �G���  �/      Some_stuffs Pv[�U  w[�U  �w[justforfun_justforfun_ [�U  ��[�U  p�[�U  p{[�U  0|[�U  ��I���  ׏/       Workout ffs �<[�U  p=[�U  �=[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0B[�U  i�`���  ��/       Meeting ffs ��Z�U  ��Z�U  @�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �Z�U  0����  ^�/       Appointment  _Z�U  �_Z�U  �`ZSome_stuffs_Some_stuffs_ �U  �cZ�U  `dZ�U   eZ�U  �eZ�U  ��t���  b�/       Workout                        justforfun_justforfun_                                       !����  T�/       Some_stuffs ��Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_ �U  `�Z�U   �Z�U  ��Z�U  `�Z�U  �$����  ��/      Birthday U  P3\�U  �3\�U  P4\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P8\�U  �����  \�/      Birthday                       This_stuffs_This_stuffs_                                     �����  �/       Some_stuffs �Z�U  PZ�U  ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Z�U  zI/���  �/       Some_stuffs ��Y�U  ��Y�U  �YThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  @�Y�U  �c����  �-�/       Workout     ��Y�U  ��Y�U  p�YSome_stuffs_Some_stuffs_ �U  ��Y�U  @�Y�U  ��Y�U  ��Y�U  �泄��  .�/       Appointment �G]�U  0H]�U  �H]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �L]�U  ���  �1�/       Workout �U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  ��ń��  �2�/      Appointment �2[�U  03[�U  �3[Some_stuffs_Some_stuffs_ �U  �5[�U  p6[�U  07[�U  �7[�U  ,)O���  �U�/      Some_stuffs 5Y�U  �5Y�U  P8Yjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  �EY�U  �$���  z}�/      Some_stuffs ��Y�U  @�Y�U  ��YSome_stuffs_Some_stuffs_ �U  ��Y�U  `�Y�U    Z�U  � Z�U  HAy���  ��/       Meeting �U   �[�U  ��[�U  @�[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��[�U  l�z���  q��/       Some_stuffs 1\�U  �1\�U  2\justforfun_justforfun_ \�U  P4\�U  �4\�U  P5\�U  6\�U  )����  ���/       Birthday    ��[�U  p�[�U  p{[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0�[�U  �鑆��  m��/       Appointment ��[�U  0�[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0�[�U  �M����  Ȩ�/      Meeting      #Z�U  �#Z�U  �$ZThis_stuffs_This_stuffs_ �U  �'Z�U  P(Z�U  )Z�U  �)Z�U  �m���  �ƀ/       Appointment �`Z�U  `aZ�U   bZSome_stuffs_Some_stuffs_ �U   eZ�U  �eZ�U  �fZ�U  0rZ�U  �g���  Xʀ/       Appointment   Z�U  � Z�U  �!ZThis_stuffs_This_stuffs_ �U  �$Z�U  p-Z�U  &Z�U  �&Z�U  r���  �ˀ/       Birthday U  �<[�U  p=[�U  �=[justforfun_justforfun_ [�U  p@[�U  �@[�U  �A[�U  0B[�U  �����  �ˀ/       Workout �U   [�U  �[�U  �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  [�U  �䢇��  O�/      Workout ffs ��Z�U  ��Z�U  0�Zjustforfun_justforfun_ _This_stuffs_This_stuffs_ �U  `�Z�U  �ޣ���  ��/       Meeting ffs �X]�U  �Y]�U  @Z]This_stuffs_This_stuffs_ �U  �\]�U   ]]�U  �]]�U  `^]�U  
s����  ��/       Workout     pf\�U  �f\�U  �g\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �k\�U  �J����  ���/       Appointment ��Y�U  `�Y�U   �YSome_stuffs_Some_stuffs_ �U  p�Y�U  0�Y�U  ��Y�U  ��Y�U  �ɼ���  ��/       Appointment 1]�U  �1]�U  @2]Some_stuffs_Some_stuffs_ �U  `4]�U  �4]�U  `5]�U  �5]�U  �|O���  ~�/      Workout     PZ�U  �Z�U  �ZThis_stuffs_This_stuffs_ �U  �Z�U  �Z�U  `Z�U   Z�U  4�ֈ��  "=�/      Birthday     �Y�U  �Y�U  0�Yjustforfun_justforfun_ Y�U  ��Y�U  ��Y�U  P�Y�U  �Y�U  �����  /A�/       Some_stuffs p�\�U  �\�U  p�\This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  ��\�U  �m���  pC�/       Appointment p�[�U  �[�U  P�[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  б[�U  ��o���  Ed�/       Appointment �<Z�U  P=Z�U  >ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  PCZ�U  Z�u���  �e�/       Some_stuffs  \Z�U  pgZ�U  �]ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �bZ�U  \q}���  �g�/      Meeting �U   �Y�U  ��Y�U  ��YSome_stuffs_Some_stuffs_ �U  P�Y�U  �Y�U  ��Y�U  ��Y�U  �v~���  h�/       Meeting      �\�U  ��\�U  @�\justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  �\�U  ��~���  h�/       Meeting     0�Z�U  ��Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0�Z�U  3�����  �h�/       Some_stuffs ��Y�U  p�Y�U  ��YThis_stuffs_This_stuffs_ �U  �Y�U  ��Y�U   �Y�U  �Y�U  T}���  v��/      Appointment                    This_stuffs_This_stuffs_                                     r�����  流/       Workout ffs  	Y�U  �	Y�U  �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `Y�U  �����  ���/       Appointment xY�U  �xY�U  �|YThis_stuffs_This_stuffs_ �U  ��Y�U  ��Y�U  p�Y�U  0�Y�U  흿���  E��/      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             $k<���  8ځ/      Appointment �0Z�U  p1Z�U  02Zjustforfun_justforfun_ _This_stuffs_This_stuffs_ �U  �7Z�U  !HT���  T��/       Appointment ��\�U   �\�U  ��\justforfun_justforfun_ _ �U  P�\�U  Щ\�U  p�\�U  0�\�U  h�ы��  q �/       Birthday U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  ��k���  �'�/      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �{���  �+�/       Some_stuffs �0Z�U  p1Z�U  02ZSome_stuffs_Some_stuffs_ �U  �4Z�U  0?Z�U  7Z�U  �7Z�U  �C���  �O�/       Workout ent 0�[�U  ��[�U  0�[This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  ��[�U  �#���  �Q�/      Some_stuffs �J\�U  PK\�U  L\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  PP\�U  �m����  nx�/       Appointment ��^�U   �^�U  ��^This_stuffs_This_stuffs_ �U  �^�U  `�^�U  �^�U  ��^�U  �����  �x�/      Workout     �Z�U  �Z�U  `ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  � Z�U  1�׎��  �Ƃ/       Appointment p�Z�U  0�Z�U  ��ZSome_stuffs_Some_stuffs_ �U  0�Z�U  � [�U  `�Z�U  ��Z�U  |����  ʂ/      Birthday U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  BXp���  ��/       Workout     �=[�U  �>[�U  p?[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pC[�U  yly���  ��/       Appointment  �Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_ �U  0�Z�U  ��Z�U  ��Z�U  p�Z�U  ,~���  -�/      Appointment p�Y�U  0�Y�U  0�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�Y�U  �c����  �/       Some_stuffs �L[�U  pM[�U  �8[Some_stuffs_Some_stuffs_ �U  p;[�U  �;[�U  �<[�U  p=[�U  �����  ��/       Appointment ��]�U  p�]�U  �]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��]�U  �����  G�/      Appointment �^�U  б^�U  P�^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P�^�U  J�����  �=�/       Some_stuffs �]�U  �]�U  0]justforfun_justforfun_ ]�U  �]�U  0]�U  �]�U  0]�U  �w����  �>�/       Some_stuffs p�\�U  0�\�U  ��\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �\�U  ������  �>�/       Workout     7Z�U  �7Z�U  P8ZThis_stuffs_This_stuffs_ �U  ;Z�U  �;Z�U  �<Z�U  P=Z�U  j�+���  1_�/       Some_stuffs ��Y�U  @�Y�U   �YSome_stuffs_Some_stuffs_ �U  ��Y�U  ��Y�U  P�Y�U  �Y�U  �<=���  �c�/       Some_stuffs 0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��X�U  �XF���  �e�/      Meeting     P*Z�U  +Z�U  �+ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �/Z�U  ځϑ��  ��/       Workout     �-Z�U  �.Z�U  0/ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  04Z�U  ��Ց��  ���/       Meeting      �X�U  ��X�U  ��XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  Y�U  Sߑ��  ��/       Birthday U  @�\�U  ��\�U  @�\justforfun_justforfun_ \�U  p�\�U  �\�U  ��\�U  P�\�U  T���  *��/       Birthday    0�]�U  ��]�U  0�]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �]�U  �����  ���/      Birthday     �Z�U  ��Z�U  `�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �Z�U  ��{���  +��/       Workout     ��\�U  `�\�U  ��\This_stuffs_This_stuffs_ �U   �\�U  ��\�U   �\�U  ��\�U  |3���  _؃/      Meeting     0MZ�U  �MZ�U  pNZSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   TZ�U  �����  ?��/       Workout     �%Y�U  �&Y�U  )YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �5Y�U  �ɰ���  F��/      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             (F���  ���/      Appointment �%Y�U  �&Y�U  )YSome_stuffs_Some_stuffs_ �U  �1Y�U  �2Y�U  5Y�U  �5Y�U  ��^���  į�/       Appointment @�\�U   �\�U  ��\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��\�U  �i���  ���/       Meeting     P�Y�U  �Y�U  ��YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �Y�U  Ox޽��  �Ў/      Meeting     �B[�U  pC[�U  0D[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0I[�U  l����  Qю/       Birthday                       Some_stuffs_Some_stuffs_                                     �2���  :Ҏ/       Appointment ��]�U  ��]�U   �]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��]�U  i����  ֎/       Workout     �m\�U   n\�U  �n\This_stuffs_This_stuffs_ �U  @q\�U   r\�U  �r\�U  @s\�U  ����  �֎/       Appointment `[�U  �[�U  �[This_stuffs_This_stuffs_ �U  �[�U  �$[�U  �[�U  P[�U  ������  �׎/       Meeting     �-Z�U  �.Z�U  0/ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  04Z�U  h����  q��/       Some_stuffs 0_[�U  �_[�U  p`[justforfun_justforfun_ [�U  Pz[�U  �z[�U  @d[�U  �d[�U  �����  ��/       Meeting ffs 0]�U  �]�U  0]This_stuffs_This_stuffs_ �U  �
]�U  0]�U  �]�U  �]�U  �����  �!�/      Some_stuffs ��X�U  ��X�U  0�Xjustforfun_justforfun_ X�U   �X�U  ��X�U  ��X�U  @�X�U  ��#���  �#�/       Workout     ��X�U  ��X�U  0�XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @�X�U  I�����  �H�/       Appointment Pu[�U  �u[�U  Pv[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p�[�U  ������  oJ�/       Birthday    �G\�U  PH\�U  �H\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �L\�U  -˿��  �N�/      Some_stuffs �Z�U  ��Z�U  p�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �Z�U  �aE���  �m�/       Workout ent ��[�U  P�[�U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P�[�U  �J���  ?o�/       Some_stuffs 0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��X�U  �*X���  �r�/      Appointment c[�U  �c[�U  N[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pR[�U  @�]���  (t�/       Birthday    p�Y�U  0�Y�U  ��YSome_stuffs_Some_stuffs_ �U  ��Y�U  ��Y�U   �Y�U  ��Y�U  ������  ���/       Birthday                       justforfun_justforfun_ _                                     �L����  ���/      Meeting      [�U  � [�U  P![This_stuffs_This_stuffs_ �U  �#[�U  p8[�U  p%[�U  0&[�U  ᱅���  쿏/       Meeting ent `5]�U  �5]�U  �6]Some_stuffs_Some_stuffs_ �U  �8]�U  `9]�U  �9]�U  �:]�U  �ʈ���  ���/       Meeting     xY�U  �xY�U  �|YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0�Y�U  �����  z�/       Meeting     0�[�U  ��[�U  p�[justforfun_justforfun_ [�U  �[�U  ��[�U  p�[�U  �[�U  �����  ]�/      Workout     �ZZ�U  @[Z�U   \ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `aZ�U  �P����  ��/       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             LM����  �W�/      Appointment ��Y�U  ��Y�U   �YThis_stuffs_This_stuffs_ �U  ��Y�U  ��Y�U   �Y�U  ��Y�U  �����  �X�/       Birthday    �Z�U  pZ�U  0	ZThis_stuffs_This_stuffs_ �U  �Z�U  �Z�U  �Z�U  @Z�U  �����  AZ�/       Meeting     �
[�U   [�U  �[justforfun_justforfun_ _ �U  �[�U  `[�U   [�U  �[�U  �i����  Æ�/       Workout     `�]�U  ��]�U  ��]Some_stuffs_Some_stuffs_ �U  ��]�U  p�]�U  ��]�U  ��]�U  t�����  ʆ�/      Meeting      YZ�U  �YZ�U  �ZZThis_stuffs_This_stuffs_ �U  �]Z�U  `^Z�U   _Z�U  �_Z�U  �B���  ��/       Meeting     ��\�U   �\�U  ��\Some_stuffs_Some_stuffs_ �U  ��\�U  @�\�U  ��\�U  @�\�U  �<���  Ъ�/       Workout ent �~Z�U  0Z�U  �Zjustforfun_justforfun_ Z�U  ��Z�U  ��Z�U  p�Z�U  0�Z�U  �����  x��/       Birthday    p�Y�U  0�Y�U  0�Yjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  p�Y�U  T$���  ��/      Birthday U   Z�U  �Z�U  �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  pZ�U  Dn����  l͐/      Appointment ��[�U  �[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��[�U  �cM���  0��/      Birthday nt ��[�U  P�[�U  �[justforfun_justforfun_ _ �U  ��[�U  P�[�U  ��[�U  P�[�U  �h����  ��/      Appointment �%Y�U  �&Y�U  )YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �5Y�U  �=����  !�/       Birthday nt  �\�U  ��\�U  `�\This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  ��\�U  
(i���  �A�/       Meeting �U  0TY�U   VY�U  @YYThis_stuffs_This_stuffs_ �U  paY�U  0bY�U  �eY�U  `fY�U  ��u���  	E�/      Meeting     PP]�U  �P]�U  PQ]Some_stuffs_Some_stuffs_ �U  �S]�U  pT]�U  �T]�U  �U]�U  +i����  �G�/       Some_stuffs 0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��X�U  �x����  �G�/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_              �����  �J�/       Some_stuffs                    Some_stuffs_Some_stuffs_                                     UM���  vp�/      Workout     EY�U  �EY�U  �HYjustforfun_justforfun_ Y�U  �PY�U  @QY�U  0TY�U   VY�U  0f ���  �p�/       Some_stuffs `�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_ �U  `�Z�U   �Z�U  ��Z�U  ��Z�U  ������  a��/       Workout     pP[�U  0Q[�U  �Q[justforfun_justforfun_ [�U  pT[�U  �T[�U  �U[�U  0V[�U  ͢���   ��/       Birthday    ��\�U   �\�U  ��\This_stuffs_This_stuffs_ �U  ��\�U  `�\�U   �\�U  ��\�U  ������  3��/      Birthday    �][�U  p^[�U  0_[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �z[�U  �^����  d��/       Appointment                    justforfun_justforfun_                                        I5���  ���/       Birthday    ��X�U  P�X�U   �XSome_stuffs_Some_stuffs_ �U   Y�U  � Y�U  �Y�U  pY�U  �@���  ���/      Some_stuffs �[�U  �[�U  `[Some_stuffs_Some_stuffs_ �U   [�U  �[�U  �[�U  �$[�U  |�v���  �	�/      Some_stuffs ��Y�U  ��Y�U   �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  1�����  ~�/       Workout     ��[�U  ��[�U  �[justforfun_justforfun_ [�U  ��[�U  P�[�U  �[�U  ��[�U  ������  ,�/      Workout     ��Y�U  ��Y�U  p�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  1�����  T�/       Meeting �U  ��Z�U  `�Z�U   �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  b]����  V�/       Some_stuffs pP[�U  0Q[�U  �Q[This_stuffs_This_stuffs_ �U  pT[�U  �T[�U  �U[�U  0V[�U  �����  Z�/       Workout     �n\�U  @o\�U  �o\justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  �t\�U  +*����  iZ�/       Appointment p?[�U  �?[�U  p@[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �D[�U  xj����  �Z�/       Appointment �%Y�U  �&Y�U  )YSome_stuffs_Some_stuffs_ �U  �1Y�U  �2Y�U  5Y�U  �5Y�U  ŗ=���  \~�/      Workout �U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  ��>���  �~�/       Appointment ��Y�U  ��Y�U   �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  ������  ϥ�/      Some_stuffs �[�U  ��[�U  P�[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �[�U  �7a���  ɒ/       Meeting      �\�U  ��\�U   �\Some_stuffs_Some_stuffs_ �U  @�\�U  ��\�U  @�\�U   �\�U  |�v���  Β/      Appointment �QZ�U  �RZ�U  �HZjustforfun_justforfun_ Z�U  �KZ�U  pLZ�U  0MZ�U  �MZ�U  �Oy���  /ϒ/       Meeting     0JZ�U  �JZ�U  �KZjustforfun_justforfun_ Z�U  pNZ�U  0OZ�U  �OZ�U  �PZ�U  @���  ���/       Meeting     0D[�U  �D[�U  �E[Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  pJ[�U  ��I���  ŝ/      Appointment p%[�U  0&[�U  �&[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p+[�U  �f����  ��/       Meeting     �_]�U  ``]�U  a]Some_stuffs_Some_stuffs_ �U  pc]�U  �c]�U  �d]�U  0e]�U  �� ���  ��/      Appointment ��Y�U  ��Y�U  p�YThis_stuffs_This_stuffs_ �U  ��Y�U  @�Y�U  ��Y�U  ��Y�U  ����  :��/       Some_stuffs 2\�U  �2\�U  P3\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  7\�U  �&y���  ��/       Appointment `�Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  E�}���  ��/      Some_stuffs �Z�U  �Z�U  �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Z�U  �����  ��/       Meeting     P�[�U  �[�U  й[justforfun_justforfun_ [�U  P�[�U  �[�U  н[�U  ��[�U  %<����  �`�/       Workout     ��[�U  P�[�U  ��[This_stuffs_This_stuffs_ �U  �[�U  ��[�U  �[�U  ��[�U  t^����  fb�/       Workout     �Z�U  PZ�U  ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Z�U  ������  �d�/       Some_stuffs �+Z�U  �,Z�U  �5ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p1Z�U  �\����  �e�/      Meeting      �\�U  ��\�U  @�\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��\�U  *]����  Ih�/       Appointment ��Z�U  ��Z�U  p�ZThis_stuffs_This_stuffs_ �U   �Z�U  ��Z�U  0�Z�U  ��Z�U  ������  dh�/       Appointment ��\�U  p�\�U  0�\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p�\�U  �tF���  ҈�/      Workout                        justforfun_justforfun_                                       ��I���  ���/       Birthday    ��\�U   �\�U  ��\Some_stuffs_Some_stuffs_ �U  ��\�U  `�\�U   �\�U  ��\�U  �`���  b��/       Birthday    @!\�U  �!\�U  p"\Some_stuffs_Some_stuffs_ �U  �$\�U  P%\�U  &\�U  �&\�U  ������  g��/      Workout     ��X�U  ��X�U  0�Xjustforfun_justforfun_ X�U   �X�U  ��X�U  ��X�U  @�X�U  @����  �۞/       Some_stuffs p�]�U  �]�U  ��]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�]�U  �����  /��/       Birthday    ��^�U  `�^�U  �^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �^�U  \����  ���/      Some_stuffs �V[�U  �W[�U  pX[This_stuffs_This_stuffs_ �U  0[[�U  �[[�U  0\[�U  �\[�U  Qv���  ��/       Birthday    ��]�U   ^�U  � ^This_stuffs_This_stuffs_ �U  �^�U  ^�U  �^�U  ^�U  �����  w(�/       Appointment @�[�U  ��[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �[�U  p�����  �)�/       Birthday U  `�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U   �Z�U  F�����  l*�/      Some_stuffs p3Z�U  04Z�U  �4ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P:Z�U  �8����  �u�/      Some_stuffs pNZ�U  0OZ�U  �OZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �UZ�U  Y����  �z�/       Some_stuffs �V[�U  �W[�U  pX[justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  �\[�U  �}���  �/      Meeting      �Z�U  ��Z�U   �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  0z  �  >ş/       Meeting ent PM\�U  �M\�U  PN\Some_stuffs_Some_stuffs_ �U  �P\�U  PQ\�U  �Q\�U  PR\�U  �++  �  �ɟ/       Workout     ��Z�U  ��Z�U  p�ZThis_stuffs_This_stuffs_ �U   �Z�U  ��Z�U  0�Z�U  ��Z�U  uO�  �  
�/      Appointment  _Z�U  �_Z�U  �`ZThis_stuffs_This_stuffs_ �U  �cZ�U  `dZ�U   eZ�U  �eZ�U  ��  �  *�/       Meeting                        This_stuffs_This_stuffs_                                     �e: �  ��/      Some_stuffs 0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��X�U  ��L �  ��/       Some_stuffs @l^�U  �l^�U  pm^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @q^�U  y�L �  ��/       Workout �U  �[�U  ��[�U  �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��[�U  r<� �  &9�/       Some_stuffs ��^�U  @�^�U  ��^Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  @�^�U  p�� �  f<�/       Meeting �U  �.[�U  p/[�U  �/[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p4[�U  ��� �  �=�/      Birthday    @�Z�U  ��Z�U  ��ZSome_stuffs_Some_stuffs_ �U  ��Z�U   �Z�U   �Z�U  ��Z�U  ��z �  a�/      Workout      �Y�U  ��Y�U  ��YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Z�U  ��| �  ya�/       Some_stuffs  |\�U  �|\�U  @}\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��\�U  ,& �  ͌�/      Workout     ��X�U  @�X�U   YThis_stuffs_This_stuffs_ �U  PY�U  Y�U   	Y�U  �	Y�U  �)� �  ��/       Meeting     ��Z�U  `�Z�U   �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `�Z�U  �J� �  歠/      Some_stuffs @�[�U   �[�U   �[Some_stuffs_Some_stuffs_ �U  @�[�U  ��[�U  ��[�U  �[�U  XN� �  筠/       Workout     &Z�U  �&Z�U  �'ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �,Z�U  }� �  ʱ�/       Some_stuffs p�Z�U  0�Z�U   �ZSome_stuffs_Some_stuffs_ �U  ��Z�U  p�Z�U  0�Z�U  ��Z�U  HQ �  ]٠/       Appointment @q]�U  �q]�U  @r]justforfun_justforfun_ _ �U  @t]�U  �t]�U  @u]�U   v]�U  0�� �  ���/       Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             Eq� �  L��/      Some_stuffs ��[�U  P�[�U  ��[Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  `�[�U  �Sh �  � �/       Appointment P�[�U  ж[�U  P�[justforfun_justforfun_ [�U  й[�U  ��[�U  �[�U  л[�U  *� �  �&�/       Appointment �e[�U   f[�U  �f[justforfun_justforfun_ [�U  @i[�U  �i[�U  @j[�U  �j[�U  �^� �  )�/       Birthday    >Z�U  pHZ�U  �?ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �DZ�U  �] �  K�/      Workout �U  ��^�U   �^�U  ��^Some_stuffs_Some_stuffs_ �U  0�^�U  ��^�U  0�^�U  ��^�U  ��� �  8n�/       Workout     Z�U  �Z�U  �Zjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  �Z�U  \<� �  �n�/       Meeting     PN\�U  �N\�U  �O\This_stuffs_This_stuffs_ �U  �Q\�U  PR\�U  S\�U  �S\�U  3� �  �p�/       Workout     й[�U  ��[�U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  п[�U  � �  .r�/      Birthday    pO[�U  �O[�U  pP[Some_stuffs_Some_stuffs_ �U  0S[�U  �S[�U  pT[�U  �T[�U  j	� �  qr�/       Meeting     ��[�U  �[�U  ��[This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ��[�U  �LG �  x��/       Some_stuffs p�[�U  0�[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p�[�U  ��� �  ���/       Workout     @i[�U  �i[�U  @j[Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  �n[�U  �� �  ���/      Meeting      {\�U  �{\�U   |\justforfun_justforfun_ \�U  @~\�U  �~\�U  @\�U  �\�U  �� �  L��/       Meeting     ��]�U  p�]�U  ��]This_stuffs_This_stuffs_ �U  ��]�U  ��]�U  �]�U  ��]�U  ��	 �  ��/       Some_stuffs ppZ�U  0qZ�U  p}ZSome_stuffs_Some_stuffs_ �U  0tZ�U  �tZ�U  puZ�U  0vZ�U  �2	 �  ��/      Some_stuffs  [�U  �[�U  �[Some_stuffs_Some_stuffs_ �U  [�U  �[�U  P[�U  [�U  !��	 �  �7�/       Workout     @i]�U  �i]�U  @j]This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  @n]�U  <�	 �  79�/      Birthday    �.[�U  p/[�U  �/[This_stuffs_This_stuffs_ �U  �2[�U  03[�U  �3[�U  p4[�U  �r0
 �  :Z�/      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �1
 �  �Z�/       Workout     ��[�U  �[�U  ��[justforfun_justforfun_ [�U  �[�U  ��[�U  P�[�U  ��[�U  ���3 �  �	�/      Some_stuffs Pu[�U  �u[�U  Pv[This_stuffs_This_stuffs_ �U  �x[�U  �y[�U  ��[�U  p�[�U  (��3 �  	�/       Workout     �rZ�U  psZ�U  0tZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �xZ�U  �}4 �  ^.�/      Birthday    `�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `�Z�U  )=�4 �  I4�/       Appointment p}Z�U  �}Z�U  �rZjustforfun_justforfun_ Z�U  puZ�U  0vZ�U  �vZ�U  pwZ�U  ���5 �  ��/       Appointment  	Y�U  �	Y�U  �YThis_stuffs_This_stuffs_ �U  �Y�U  `Y�U  �Y�U  `Y�U  ���5 �  ���/      Some_stuffs  YZ�U  �YZ�U  �ZZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �_Z�U  }H6 �  ߣ�/      Appointment 0S[�U  �S[�U  pT[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0Y[�U  B�_6 �  詭/       Some_stuffs P![�U  "[�U  �"[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0'[�U  ��b6 �  ���/       Appointment @�Z�U  ��Z�U  �ZSome_stuffs_Some_stuffs_ �U  p�Z�U  ��Z�U  ��Z�U  p�Z�U  ��6 �  �ѭ/      Birthday    0MZ�U  �MZ�U  pNZjustforfun_justforfun_ Z�U  �\Z�U   ]Z�U  @SZ�U   TZ�U  <��7 �  w��/      Workout     p�Y�U  0�Y�U  0�YSome_stuffs_Some_stuffs_ �U   �Y�U  ��Y�U  ��Y�U  p�Y�U  "&�7 �  ��/       Birthday    PF\�U  G\�U  �G\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  PK\�U  A��7 �  ���/       Appointment �[�U  ��[�U  p�[justforfun_justforfun_ [�U  ��[�U  �[�U  ��[�U  P�[�U  O�8 �  A�/      Birthday    ��]�U  �]�U  ��]Some_stuffs_Some_stuffs_ �U  �^�U  ^�U  �^�U  ^�U  ʌ8 �  M�/       Some_stuffs �Y�U  `Y�U  �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �&Y�U  o!8 �  
�/       Some_stuffs �`Z�U  `aZ�U   bZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0rZ�U  8�!8 �  �/       Some_stuffs �jZ�U  pkZ�U  0lZSome_stuffs_Some_stuffs_ �U  �nZ�U  �oZ�U  ppZ�U  0qZ�U  ��!8 �  %�/       Birthday    ��Y�U  ��Y�U  P�YSome_stuffs_Some_stuffs_ �U  �Y�U  ��Y�U  0�Y�U  ��Y�U   ��8 �  @E�/       Some_stuffs @l\�U  �l\�U  �m\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   r\�U  )��8 �  �F�/       Birthday    ��[�U  ��[�U  @�[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @�[�U  ��D9 �  �g�/       Some_stuffs �Z�U  �Z�U  �ZSome_stuffs_Some_stuffs_ �U  0	Z�U  �	Z�U  p
Z�U  0Z�U  �c9 �  ]o�/      Birthday    ��Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `�Z�U  �=�9 �  I��/      Meeting                        Some_stuffs_Some_stuffs_                                     �~: �  ѷ�/      Birthday nt ��Y�U  �Y�U  ��Yjustforfun_justforfun_ _This_stuffs_This_stuffs_ �U  @�Y�U  ɤ�: �  M��/       Workout  U  �J^�U  PK^�U  �K^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �O^�U  Z�: �  缮/       Meeting ffs ��^�U  `�^�U  ��^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��^�U  ��; �  �߮/      Birthday                       Some_stuffs_Some_stuffs_                                     �E; �  �/       Some_stuffs @�\�U  ��\�U  @�\justforfun_justforfun_ \�U  ��\�U  P�\�U  Л\�U  ��\�U  �"; �   �/       Appointment �[�U  p�[�U  0�[justforfun_justforfun_ [�U  �[�U  p�[�U  0�[�U  �[�U  4��; �  ��/      Meeting �U  ��Z�U  ��Z�U  @�ZSome_stuffs_Some_stuffs_ �U   �Z�U  ��Z�U  ��Z�U   �Z�U   9J< �  �-�/       Meeting     5Y�U  �5Y�U  P8YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �EY�U  �O< �  �.�/      Workout     �eY�U  `fY�U  �iYjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  �xY�U  ���< �  /U�/       Some_stuffs ��Z�U  p�Z�U  0�Zjustforfun_justforfun_ Z�U  ��Z�U  0�Z�U  ��Z�U  ��Z�U  �t�< �  �V�/      Some_stuffs ��[�U  ��[�U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��[�U  @��= �  h��/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ���= �  /      Workout     �a[�U  0b[�U  Pz[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @g[�U  ��$> �  ��/       Meeting  nt ��]�U  @�]�U  ��]This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  @�]�U  �0(> �  ���/      Birthday    �|[�U  p}[�U  0~[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��[�U  !�9? �  ��/       Appointment �Z�U  �Z�U  PZjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  �Z�U  �CQ? �  	��/      Workout     N[�U  �N[�U  pO[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �S[�U  ���? �  :�/      Birthday fs 0�[�U  ��[�U  0�[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  Ь[�U  ��? �  ��/       Birthday    @�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_ �U  ��Z�U  `�Z�U   �Z�U  ��Z�U  ��z@ �  7@�/       Workout     �[�U  ��[�U  ��[justforfun_justforfun_ [�U  �[�U  ��[�U  ��[�U  �[�U  J~@ �  A�/      Appointment ��Y�U  @�Y�U  ��YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  	�A �  �f�/       Birthday    �\�U  ��\�U  �\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��\�U  �A �  j�/       Some_stuffs `\�U  �\�U  `\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `\�U  hX�A �  щ�/       Appointment ��Y�U  `�Y�U   �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  A�A �  ��/       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �q�A �  D��/       Meeting     �Z�U  ��Z�U   �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Z�U  x>B �  ճ�/       Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             sEB �  ���/       Some_stuffs  �Y�U  ЕY�U   �Yjustforfun_justforfun_ Y�U  ��Y�U  p�Y�U  ��Y�U  ��Y�U  R*IB �  ���/       Some_stuffs  ]\�U  �]\�U  P^\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �b\�U  U�LB �  v��/      Birthday    �eY�U  `fY�U  �iYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �xY�U  H`�B �  }۰/       Some_stuffs �[�U  p�[�U  0�[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��[�U  �^�B �  �ް/      Birthday    0 ]�U  � ]�U  0]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p]�U  [�bC �  ���/       Appointment s[�U  �s[�U  t[Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  Px[�U  �eC �  `��/       Appointment ��Y�U  ��Y�U   �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  ��tC �  K�/       Appointment �Z�U  pZ�U  0	ZThis_stuffs_This_stuffs_ �U  �Z�U  �Z�U  �Z�U  @Z�U  ���C �  �/      Some_stuffs p�[�U  0�[�U  ��[Some_stuffs_Some_stuffs_ �U  p�[�U  �[�U  P�[�U  �[�U  ͂D �  (�/      Meeting     P^\�U  �^\�U  @�\This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  �c\�U  H�D �  )�/       Birthday    p�Z�U  0�Z�U  ��ZSome_stuffs_Some_stuffs_ �U  ��Z�U  ��Z�U  p�Z�U  ��Z�U  ,#5E �  v�/      Some_stuffs �!Z�U  @"Z�U   #ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P(Z�U  QGGE �  �z�/       Meeting �U  �/^�U   0^�U  �0^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   5^�U  ��o �  �K�/       Workout      �]�U  ��]�U   �]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��]�U  �/�o �  �P�/       Meeting     7Z�U  �7Z�U  P8Zjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  P=Z�U  �J�o �  �Q�/      Meeting ent @�[�U  ��[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �[�U  `^p �  �p�/       Some_stuffs `�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_ �U  `[�U   [�U  �[�U  `[�U  #�p �  Tq�/       Birthday     �Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_ �U  ��Z�U  ` [�U  `[�U   [�U  �*p �  lu�/       Workout �U  ��[�U  ��[�U  �[Some_stuffs_Some_stuffs_ �U  ��[�U  P�[�U  �[�U  ��[�U  ͋3p �  �w�/      Workout     ��Z�U  ��Z�U  0�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0�Z�U  :ȼp �  Ӛ�/       Some_stuffs �Z�U  pZ�U  0	ZThis_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  @Z�U  )��p �  	��/       Some_stuffs  �^�U  ��^�U   �^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��^�U  (��p �  )��/       Appointment �?]�U  `@]�U   A]Some_stuffs_Some_stuffs_ �U  �C]�U  D]�U  �D]�U  E]�U  5Oq �  b��/      Birthday    �[�U  �[�U   [This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p8[�U  ��Oq �  d��/       Birthday    p�Z�U  0�Z�U  ��ZThis_stuffs_This_stuffs_ �U  ��Z�U  ��Z�U  p�Z�U  ��Z�U  �~�q �  �/       Workout      	Y�U  �	Y�U  �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `Y�U  ���q �  ��/       Appointment �	\�U  �
\�U   \justforfun_justforfun_ \�U  �\�U  p\�U  0\�U  �\�U  ���q �  �/       Workout     ��X�U  @�X�U   YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �	Y�U  �I�q �  �/      Meeting     EY�U  �EY�U  �HYThis_stuffs_This_stuffs_ �U  �PY�U  @QY�U  0TY�U   VY�U  ��r �  $�/       Appointment  ;]�U  �;]�U  �<]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `@]�U  D+�r �  ��/      Some_stuffs   Z�U  � Z�U  �!ZThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  �&Z�U  R�#s �  28�/       Some_stuffs P�^�U  Ќ^�U  ��^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0�^�U  ��)s �  �9�/       Birthday    ��Y�U  ��Y�U   �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  ��/s �  S;�/      Appointment                    This_stuffs_This_stuffs_                                     �o�s �  X_�/       Birthday    �Z�U  pZ�U  0	ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @Z�U  ���s �  �_�/       Meeting      �]�U  ��]�U  0�]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �]�U  ��_t �  1��/      Birthday    @�Z�U   �Z�U  ��Zjustforfun_justforfun_ Z�U  ��Z�U   �Z�U  ��Z�U  ��Z�U   ��t �   ��/       Meeting     �Z�U  pZ�U  0	ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @Z�U  q��t �  &��/       Some_stuffs p�]�U  �]�U  p�]This_stuffs_This_stuffs_ �U  ��]�U  @�]�U  0�]�U  ��]�U  �t �  `��/       Birthday    @�\�U  P�\�U  ��\justforfun_justforfun_ \�U  ��\�U  @�\�U  ��\�U  ��\�U  ���t �  G��/      Appointment  �Z�U  ��Z�U   �Zjustforfun_justforfun_ _This_stuffs_This_stuffs_ �U  ��Z�U  ��vu �  �н/       Meeting ffs �'[�U  p([�U  0)[This_stuffs_This_stuffs_ �U  0,[�U  �,[�U  p-[�U  �-[�U  h߄u �  1Խ/       Workout     ��Y�U  ��Y�U  p�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  ]t�u �  �׽/      Some_stuffs �\�U  p\�U  �\justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  �!\�U  ZRv �  g��/       Workout ffs P3\�U  �3\�U  P4\justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  P8\�U  �cv �  0��/       Some_stuffs  _Z�U  �_Z�U  �`ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �eZ�U  ��v �  ���/      Some_stuffs ��X�U  ��X�U  0�XThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @�X�U  ��v �  ���/       Workout ffs �<[�U  p=[�U  �=[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0B[�U  ��v �  ��/       Appointment ��Y�U  `�Y�U    ZThis_stuffs_This_stuffs_ �U   Z�U  �Z�U  �Z�U   Z�U  R��v �  � �/       Meeting     PS^�U  �S^�U  �T^justforfun_justforfun_ _ his_stuffs_This_stuffs_ �U  PX^�U  ���v �  �"�/      Appointment �[�U  ��[�U  P�[justforfun_justforfun_ [�U   �[�U  ��[�U  @�[�U  ��[�U  �v �  U#�/       Appointment �+Z�U  �,Z�U  �5ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p1Z�U  ��Ow �  �I�/      Birthday U  `�Z�U   �Z�U  ��Zjustforfun_justforfun_ [�U  `[�U   [�U  �[�U  `[�U  �Sw �  �J�/       Birthday    7Z�U  �7Z�U  P8ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P=Z�U  ص�w �  �q�/       Appointment ��Z�U  ��Z�U  p�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0�Z�U  ��zx �  +��/       Some_stuffs ��\�U  `�\�U  ��\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @�\�U  �
�x �  䚾/       Meeting ent �Z�U  @Z�U  PZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  PZ�U  bh
y �  ���/       Appointment г[�U  ��[�U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �[�U  i�y �  ���/       Meeting ffs �Z�U  ��Z�U  p�ZSome_stuffs_Some_stuffs_ �U  p�Z�U  0�Z�U  ��Z�U  ��Z�U  ;�y �  ���/       Some_stuffs  �]�U  ��]�U  `�]Some_stuffs_Some_stuffs_ �U  ��]�U   �]�U  ��]�U   �]�U  ��y �  ���/       Some_stuffs P�Y�U  �Y�U  ��YThis_stuffs_This_stuffs_ �U   �Y�U  ��Y�U  ��Y�U  ��Y�U  щ�y �  B�/       Appointment `\�U   \�U  �\Some_stuffs_Some_stuffs_ �U  0\�U  �\�U  �\�U  p\�U  l��y �  �/      Workout     ��Y�U  @�Y�U  ��YThis_stuffs_This_stuffs_ �U  ��Y�U  ��Y�U  `�Y�U   �Y�U  Y7=z �  �	�/       Birthday    �[�U  ��[�U  ��[justforfun_justforfun_ [�U  ��[�U  P�[�U  �[�U  ��[�U  ��Dz �  z�/      Workout                        justforfun_justforfun_                                       3Qz �  ��/       Appointment ��Y�U  ��Y�U  `�YThis_stuffs_This_stuffs_ �U  ��Y�U  ��Y�U  p�Y�U  0�Y�U  �Vz �  
�/       Workout     `�]�U  �]�U  ��]Some_stuffs_Some_stuffs_ �U  � ^�U  ^�U  �^�U  ^�U  �Xz �  ��/       Appointment @�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @�Z�U  ��Yz �  ��/       Meeting     ��\�U  ��\�U  0�\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @�\�U  ��z �  A/�/       Some_stuffs  �Z�U  �Z�U  `�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  Z�z �  G5�/       Appointment pT[�U  �T[�U  �U[justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  pZ[�U  ��z �  D7�/      Some_stuffs �Z�U  PZ�U  ZSome_stuffs_Some_stuffs_ �U  `Z�U   Z�U  �Z�U  �Z�U  �m{ �  OW�/       Birthday    ��\�U  p�\�U  �\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �\�U  ��q{ �  xX�/       Birthday U  ��X�U  @�X�U   YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �	Y�U  ��~{ �  �[�/       Birthday    �gZ�U  phZ�U  0iZThis_stuffs_This_stuffs_ �U  0lZ�U  �lZ�U  pmZ�U  0nZ�U  �^| �  邿/      Workout     ��[�U  0�[�U  �[justforfun_justforfun_ [�U  p�[�U  0�[�U  �[�U  p�[�U  ):| �  i��/       Appointment ��^�U  @�^�U  ��^This_stuffs_This_stuffs_ �U  ��^�U  @�^�U  ��^�U  p�^�U  �N�| �  ���/       Meeting     ��[�U  ��[�U   �[justforfun_justforfun_ _ �U  ��[�U  @�[�U  ��[�U  ��[�U   @} �  �ο/      Appointment ��[�U  P�[�U  ��[This_stuffs_This_stuffs_ �U  ��[�U  �[�U  ��[�U  P�[�U  0fG} �  �п/       Appointment pc]�U  �c]�U  �d]Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  �h]�U  ��} �  ���/      Workout     PAZ�U  �AZ�U  �BZSome_stuffs_Some_stuffs_ �U  �EZ�U  PFZ�U  GZ�U  �GZ�U  Ćd~ �  ��/      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_              � �  �C�/       Meeting �U  P�Y�U  �Y�U  ��YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  �r �  �D�/       Some_stuffs ��Z�U  0�Z�U  �ZThis_stuffs_This_stuffs_ �U  ��Z�U  0�Z�U  �Z�U  ��Z�U  Y� �  �H�/       Appointment P�Y�U  �Y�U  ��YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  6$ �  �I�/      Meeting      �\�U  ��\�U   �\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �\�U  q�� �  �j�/       Workout     P�[�U  п[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��[�U  <�� �  7l�/      Appointment @j[�U  �j[�U  @k[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �o[�U  �L� �  vp�/       Birthday    �Z�U  �Z�U  �ZSome_stuffs_Some_stuffs_ �U  0	Z�U  �	Z�U  p
Z�U  0Z�U  h�K� �  q��/       Workout     9^�U  �9^�U  p:^justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  P>^�U  �y΀ �  ��/       Birthday    `�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_ �U   �Z�U  ��Z�U  `�Z�U  ��Z�U  L�Ԁ �  ���/      Meeting     �L[�U  pM[�U  �8[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p=[�U  �*b� �  ���/      Workout     P^\�U  �^\�U  @�\This_stuffs_This_stuffs_ �U  �a\�U  �b\�U  pc\�U  �c\�U  y�e� �  ���/       Birthday    ��Z�U  ��Z�U  @�ZThis_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  ��Z�U  ��[(�  �T
 /      Birthday    ��Y�U  @�Y�U  ��YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  i8_(�  �U
 /       Appointment  �Y�U  ��Y�U  ��YThis_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  ЕY�U  ���(�  :y
 /      Workout     �Z�U  �Z�U  �Zjustforfun_justforfun_ Z�U  0	Z�U  �	Z�U  p
Z�U  0Z�U  [��(�  '}
 /       Appointment ��Z�U  @�Z�U   �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Z�U  hl�(�  Q~
 /       Workout     ��Y�U  ��Y�U  p�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  �� )�  8
 /       Meeting      	Y�U  �	Y�U  �YSome_stuffs_Some_stuffs_ �U  �Y�U  `Y�U  �Y�U  `Y�U  �[�)�  ֟
 /       Birthday fs  �]�U  ��]�U   �]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �]�U  ㍆)�  l�
 /       Some_stuffs ��]�U   �]�U  ��]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P�]�U  �<�)�  "�
 /       Some_stuffs @�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  @�Z�U  �D�)�  ��
 /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �*�  ��
 /       Some_stuffs �2^�U  �3^�U  `4^This_stuffs_This_stuffs_ �U  �6^�U  07^�U  �7^�U  P8^�U  ��%*�  <�
 /      Some_stuffs EY�U  �EY�U  �HYjustforfun_justforfun_ Y�U  �PY�U  @QY�U  0TY�U   VY�U  �e4*�  ��
 /       Appointment ��Y�U  ��Y�U  p�YThis_stuffs_This_stuffs_ �U  ��Y�U  @�Y�U  ��Y�U  ��Y�U  ]R�*�  k�
 /      Some_stuffs ��Y�U  ��Y�U  p�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  Hz�*�  ��
 /       Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             Jٽ*�  �
 /       Appointment �Y�U  `Y�U  �YThis_stuffs_This_stuffs_ �U  �"Y�U  `#Y�U  �%Y�U  �&Y�U  z#W+�  [ /       Appointment �o\�U  �p\�U  @q\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   v\�U  �#W+�  [ /      Birthday    EY�U  �EY�U  �HYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   VY�U  F[+�  j /       Workout �U  @\�U  �\�U  @�\Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   �\�U  c+�  j /       Meeting �U  �(\�U  �)\�U  P*\Some_stuffs_Some_stuffs_ �U  �,\�U  P-\�U  .\�U  �.\�U  �k+�  � /       Appointment �%Y�U  �&Y�U  )YThis_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  �5Y�U  ���+�  �B /       Appointment ��\�U  `�\�U  ��\justforfun_justforfun_ \�U   �\�U  ��\�U  `�\�U  ��\�U  a~,�  �D /       Meeting     ��[�U  �[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��[�U  ��{,�  Oc /      Meeting     ��X�U  ��X�U  0�XSome_stuffs_Some_stuffs_ �U   �X�U  ��X�U  ��X�U  @�X�U  �Y-�  � /       Some_stuffs  �\�U  ��\�U  `�\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `�\�U  �-�  �� /       Workout      �]�U  ��]�U  0�]justforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U  ��]�U  mu"-�  � /       Workout     P^�U  �^�U  ��^justforfun_justforfun_ _ �U  ��^�U  @�^�U  ��^�U  @�^�U  �+-�  $� /       Some_stuffs  �Y�U  �Y�U  0�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Y�U  
O+-�  5� /       Birthday    �2[�U  03[�U  �3[Some_stuffs_Some_stuffs_ �U  �5[�U  p6[�U  07[�U  �7[�U  ��0-�  �� /      Workout      �Y�U  ��Y�U  ��Yjustforfun_justforfun_ Y�U  P�Y�U  �Y�U  ��Y�U  ��Y�U  Ľ�-�  � /      Some_stuffs ��Y�U  @�Y�U   �YSome_stuffs_Some_stuffs_ �U  ��Y�U  ��Y�U  P�Y�U  �Y�U  (6K.�  �� /       Some_stuffs  �Y�U  �Y�U  0�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Y�U  'X.�  9� /      Some_stuffs ��Z�U   �Z�U   �ZSome_stuffs_Some_stuffs_ �U  `�Z�U   �Z�U  ��Z�U  `�Z�U  L0Y.�  }� /       Appointment  �Z�U  ��Z�U  `�ZThis_stuffs_This_stuffs_ �U  ��Z�U  ��Z�U  `�Z�U   �Z�U  }�Y.�  �� /       Appointment ;Z�U  �;Z�U  �<Zjustforfun_justforfun_ Z�U  �?Z�U  �@Z�U  PAZ�U  �AZ�U  Z.�  �� /       Workout     ��X�U  @�X�U   YThis_stuffs_This_stuffs_ �U  PY�U  Y�U   	Y�U  �	Y�U  Qp\.�  R� /       Meeting �U  EY�U  �EY�U  �HYSome_stuffs_Some_stuffs_ �U  �PY�U  @QY�U  0TY�U   VY�U  q/�.�  � /       Some_stuffs  [�U  �[�U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  [�U  ���.�  ) /      Appointment �Z�U  @Z�U  PZSome_stuffs_Some_stuffs_ �U  PZ�U  �Z�U  �Z�U  PZ�U  \ʁ/�  k) /      Meeting �U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  ��0�  �M /      Meeting     ��Z�U  p�Z�U  0�ZSome_stuffs_Some_stuffs_ �U  ��Z�U  0�Z�U  �Z�U  ��Z�U  �9'0�  �S /       Appointment ��Y�U  ��Y�U  �YSome_stuffs_Some_stuffs_ �U  `�Y�U   �Y�U  ��Y�U  `�Y�U  �s�0�  Wt /       Appointment P�^�U  й^�U  P�^justforfun_justforfun_ ^�U  P�^�U  �^�U  ��^�U  �^�U  �g�0�  �u /      Workout      �Y�U  ��Y�U  ��YThis_stuffs_This_stuffs_ �U  �Z�U  `Z�U   Z�U  �Z�U  ��0�  w /       Workout     �[�U  [�U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  #[�U  ��O1�  �� /       Appointment PT\�U  �T\�U  PU\justforfun_justforfun_ \�U  �W\�U  PX\�U  Y\�U  �Y\�U  ��`1�  � /       Appointment 7Z�U  �7Z�U  P8ZThis_stuffs_This_stuffs_ �U  ;Z�U  �;Z�U  �<Z�U  P=Z�U  \��1�  �� /      Birthday     	Y�U  �	Y�U  �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `Y�U  ��2�  9� /      Meeting ent �eY�U  `fY�U  �iYjustforfun_justforfun_ _ �U  �sY�U  `tY�U  xY�U  �xY�U  ���2�  �� /       Workout     �^]�U  `_]�U  �_]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �c]�U  1_3�  ^ /       Some_stuffs  �Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_ �U  0�Z�U  ��Z�U  ��Z�U  p�Z�U  �*3�   /      Workout     ��Y�U  p�Y�U  ��YThis_stuffs_This_stuffs_ �U  �Y�U  ��Y�U   �Y�U  �Y�U  �Ҩ3�  �9 /       Birthday    �Z�U  @Z�U  PZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  PZ�U  I�3�  �9 /       Some_stuffs �\�U  p\�U  �\Some_stuffs_Some_stuffs_ �U  0\�U  �\�U  p\�U  �\�U  �ҷ3�  e= /       Birthday    0]�U  �]�U  p]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p]�U  {�3�  �> /       Some_stuffs  eZ�U  �eZ�U  �fZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  pkZ�U  �jS4�  :e /       Meeting      �Y�U  ��Y�U  ��Yjustforfun_justforfun_ Y�U  ��Y�U  ��Y�U  �Y�U  ��Y�U  ,O�4�  �� /      Some_stuffs `�Z�U   �Z�U  оZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Z�U  9q�4�  s� /       Meeting     0�[�U  �[�U  p�[Some_stuffs_Some_stuffs_ �U  0�[�U  ��[�U  0�[�U  ��[�U  +�x5�  I� /       Workout     �/\�U  P0\�U  1\Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  �4\�U  �	5�  � /       Workout �U  �QZ�U  �RZ�U  �HZjustforfun_justforfun_ Z�U  �KZ�U  pLZ�U  0MZ�U  �MZ�U  Ъ�5�  � /       Meeting �U  EY�U  �EY�U  �HYSome_stuffs_Some_stuffs_ �U  �PY�U  @QY�U  0TY�U   VY�U  ~��5�  � /      Appointment 5Y�U  �5Y�U  P8YSome_stuffs_Some_stuffs_ �U  @?Y�U  AY�U  EY�U  �EY�U  c�6�  |� /       Appointment �PY�U  @QY�U  0TYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0bY�U  �w6�  �� /       Workout     p�Z�U  0�Z�U  ��ZSome_stuffs_Some_stuffs_ �U  ��Z�U  ��Z�U  p�Z�U  ��Z�U  ��6�  �� /       Appointment 0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��X�U  �6�  �� /       Birthday    0	Z�U  �	Z�U  p
Zjustforfun_justforfun_ Z�U  �Z�U  @Z�U  PZ�U  Z�U  f�!6�  �� /      Workout �U  �U[�U  0V[�U  �V[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �[[�U  RA�6�  �� /       Appointment �]�U   ]�U  �]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �!]�U  lG�6�  5� /      Some_stuffs                    This_stuffs_This_stuffs_                                     Q@�6�  R  /       Workout     ��[�U  P�[�U  �[This_stuffs_This_stuffs_ �U  ��[�U  `�[�U  �\�U  P\�U  0�W7�  �* /       Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ���7�  �J /       Some_stuffs  	Y�U  �	Y�U  �YThis_stuffs_This_stuffs_ �U  �Y�U  `Y�U  �Y�U  `Y�U  r��7�  FM /       Workout     �[�U  0�[�U  ��[Some_stuffs_Some_stuffs_ �U  p�[�U  0�[�U  ��[�U  0�[�U  �]�7�  �N /      Some_stuffs 0�Z�U  ��Z�U  @�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �Z�U  ���7�  R /       Workout     P�Y�U  �Y�U  ��YSome_stuffs_Some_stuffs_ �U   �Y�U  ��Y�U  ��Y�U  ��Y�U  8Gf8�  3p /       Appointment P�Y�U  �Y�U  ��Yjustforfun_justforfun_ Y�U   �Y�U  ��Y�U  ��Y�U  ��Y�U  �Yp8�  �r /      Meeting     �6\�U  7\�U  �7\This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  P<\�U  j��8�  �x /       Meeting ent ��Y�U  ��Y�U  p�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  ��9�  Ě /       Meeting ffs p	]�U  0
]�U  �
]justforfun_justforfun_ ]�U  0]�U  �]�U  p]�U  �]�U  I�9�  �� /       Workout     0\�U  �\�U  0\justforfun_justforfun_ \�U  0\�U  �\�U  �\�U  0\�U  �O9�  � /       Appointment �\�U  ��\�U  ��\Some_stuffs_Some_stuffs_ �U   �\�U  ��\�U  ��\�U  `�\�U  ��9�  ^� /      Meeting     �[�U  `[�U   [This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  �[�U   �9�  4� /       Meeting     �[�U  ��[�U  �[Some_stuffs_Some_stuffs_ �U  ��[�U  ��[�U  �[�U  ��[�U  T<:�  v� /      Some_stuffs �[�U  P[�U  �[This_stuffs_This_stuffs_ �U  �[�U  [�U  �[�U  �[�U  ��c�  A� /       Some_stuffs �w[�U  Px[�U  �x[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p}[�U  4u�c�  "� /      Appointment �[�U  p�[�U  0�[justforfun_justforfun_ [�U  ��[�U  p�[�U  0�[�U  ��[�U  \7�d�  �� /      Workout �U  �Z�U  PZ�U  Zjustforfun_justforfun_ Z�U  `Z�U   Z�U  �Z�U  �Z�U  ��e�  �� /       Some_stuffs  �Z�U  ��Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �Z�U  e�e�  @� /      Appointment 0[[�U  �[[�U  0\[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �`[�U  ��;e�  p� /       Workout     P^�U  �^�U  P^Some_stuffs_Some_stuffs_ �U  p^�U  �^�U  p^�U  0^�U  �=e�  �� /       Some_stuffs `�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_ �U   �Z�U  ��Z�U  `�Z�U  ��Z�U  �)�e�  s /      Appointment �EZ�U  PFZ�U  GZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �JZ�U  ��lf�  }8 /      Birthday U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��X�U  :�f�  W /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ���f�  e\ /       Appointment ��Z�U  ��Z�U  p�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  ܇g�  �~ /      Appointment ��X�U  @�X�U   YSome_stuffs_Some_stuffs_ �U  PY�U  Y�U   	Y�U  �	Y�U  �w�g�  �� /       Some_stuffs �V[�U  �W[�U  pX[This_stuffs_This_stuffs_ �U  0[[�U  �[[�U  0\[�U  �\[�U  ���g�  �� /       Some_stuffs 0�\�U  ��\�U  0 ]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0]�U  {�g�  [� /       Appointment @�[�U  ��[�U  @�[This_stuffs_This_stuffs_ �U  ��[�U  @�[�U   �[�U  ��[�U  A�h�  ȥ /       Birthday U  ��Y�U  ��Y�U  �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `�Y�U  �@h�  �� /      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �.,h�  � /       Appointment �<Z�U  P=Z�U  >ZThis_stuffs_This_stuffs_ �U  PAZ�U  �AZ�U  �BZ�U  PCZ�U  �^�h�  �� /       Meeting     pd\�U  �d\�U  pe\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �i\�U  ��h�  � /       Birthday     _Z�U  �_Z�U  �`ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �eZ�U  cv�h�  �� /       Meeting �U  �^�U  ��^�U  @�^justforfun_justforfun_ ^�U  ��^�U   �^�U  ��^�U   �^�U  �C�h�  2� /      Meeting     �]�U  0]�U  �]Some_stuffs_Some_stuffs_ �U  p]�U  0]�U  �]�U  0]�U  �Ui�  � /       Meeting     ��[�U  p�[�U  0�[justforfun_justforfun_ [�U  0�[�U  ��[�U  p�[�U  0�[�U  3�Vi�  ~� /       Workout ffs оZ�U  P�Z�U  0�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Z�U  �ei�  %� /       Some_stuffs 5Y�U  �5Y�U  P8YSome_stuffs_Some_stuffs_ �U  @?Y�U  AY�U  EY�U  �EY�U  <Ifi�  w� /      Appointment 0lZ�U  �lZ�U  pmZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �}Z�U  L�gi�  �� /       Workout �U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��X�U  ���i�  g /      Workout ffs �Z�U  �Z�U  PZSome_stuffs_Some_stuffs_ �U  Z�U  �Z�U  �Z�U  �Z�U  �K�i�  � /       Workout ent �F]�U  0G]�U  �G]Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  �K]�U  @��i�  � /       Some_stuffs ppZ�U  0qZ�U  p}Zjustforfun_justforfun_ Z�U  0tZ�U  �tZ�U  puZ�U  0vZ�U  ���i�  9! /       Meeting                        This_stuffs_This_stuffs_                                     D<�j�  (D /       Workout ffs �7\�U  P8\�U  �8\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �=\�U  K��j�  }D /       Workout ffs �Z�U  �Z�U  `ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �%Z�U  ڥ�j�  �G /       Birthday U  @�\�U  P�\�U  ��\Some_stuffs_Some_stuffs_ �U  ��\�U  @�\�U  ��\�U  ��\�U  �؏j�  �G /       Some_stuffs 01[�U  �1[�U  �2[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p6[�U  ŉ�j�  �I /      Workout     5Y�U  �5Y�U  P8YSome_stuffs_Some_stuffs_ �U  @?Y�U  AY�U  EY�U  �EY�U  ��,k�  �o /      Meeting     &Z�U  �&Z�U  �'ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �,Z�U  ��2k�  Pq /       Some_stuffs �Z�U  ��Z�U   �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Z�U  X��k�  � /       Birthday    EY�U  �EY�U  �HYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   VY�U  Bz�k�  � /       Appointment �g^�U  @h^�U  �h^Some_stuffs_Some_stuffs_ �U  �j^�U  �k^�U  @l^�U  �l^�U  ���k�  �� /      Appointment 0�Z�U  �Z�U  p�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Z�U  ��@l�  �� /       Birthday    `�Z�U  ��Z�U  `�Zjustforfun_justforfun_ Z�U   �Z�U  ��Z�U  `�Z�U  ��Z�U  t�Hl�  �� /      Some_stuffs p�Y�U  0�Y�U  0�YSome_stuffs_Some_stuffs_ �U   �Y�U  ��Y�U  ��Y�U  p�Y�U  �M�l�  t� /      Some_stuffs �a[�U  0b[�U  Pz[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @g[�U  X�l�  �� /       Workout     �Z�U  ��Z�U  p�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  ��l�  ,� /       Some_stuffs �Z�U  �Z�U  `ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  � Z�U  1 �m�  � /       Workout     `�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Z�U  r	�m�  F /       Appointment �[�U  ��[�U  ��[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��[�U  �Ԏm�  � /      Meeting     ��[�U  ��[�U  @�[This_stuffs_This_stuffs_ �U  ��[�U  ��[�U  �[�U  ��[�U   i
n�  �+ /       Meeting     ��X�U  P�X�U   �XThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  pY�U  E�n�  l, /      Workout �U  0K[�U  �K[�U  c[justforfun_justforfun_ [�U  pO[�U  �O[�U  pP[�U  0Q[�U  �~#n�  2 /       Birthday    PT\�U  �T\�U  PU\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Y\�U  �3)n�  �3 /       Birthday    DZ�U  �DZ�U  �EZSome_stuffs_Some_stuffs_ �U  �QZ�U  �RZ�U  �HZ�U  �IZ�U  x#�n�  [X /       Some_stuffs ��Z�U  0�Z�U  �Zjustforfun_justforfun_ Z�U  �Z�U  p�Z�U  ��Z�U  ��Z�U  �Go�  �| /       Workout     p�Y�U  0�Y�U  0�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p�Y�U  �&Vo�  �� /       Meeting     �Z�U  p�Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  ��]o�  r� /      Birthday    ��Z�U  0�Z�U  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  K_�o�  ݠ /       Some_stuffs  �]�U  ��]�U   �]justforfun_justforfun_ ]�U   �]�U  ��]�U   �]�U  ��]�U  ���o�  k� /       Appointment �9]�U  �:]�U   ;]Some_stuffs_Some_stuffs_ �U  �=]�U   >]�U  �>]�U  `?]�U  x��o�  �� /       Workout ent P[�U  [�U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  "[�U  ��o�  �� /      Appointment p�Y�U  0�Y�U  0�YThis_stuffs_This_stuffs_ �U   �Y�U  ��Y�U  ��Y�U  p�Y�U  :op�  s� /       Some_stuffs ��[�U  p�[�U  0�[Some_stuffs_Some_stuffs_ �U  ��[�U  0�[�U  ��[�U  p�[�U  YH�p�  '� /       Workout       Z�U  � Z�U  �!ZSome_stuffs_Some_stuffs_ �U  �$Z�U  p-Z�U  &Z�U  �&Z�U  ��p�  '� /      Meeting �U  p�Z�U  0�Z�U  ��ZThis_stuffs_This_stuffs_ �U  ��Z�U  ��Z�U  p�Z�U  ��Z�U  �'�p�  +� /       Some_stuffs 0_[�U  �_[�U  p`[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �d[�U  �cq�  �� /       Meeting     �+Z�U  �,Z�U  �5ZThis_stuffs_This_stuffs_ �U  0/Z�U  �/Z�U  �0Z�U  p1Z�U  |$q�  �� /       Birthday nt @}\�U  �}\�U  @~\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �\�U  �Zq�  � /       Workout �U  p`[�U  �`[�U  �a[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   f[�U  �}q�  �� /      Workout     ��Y�U  ��Y�U   �YThis_stuffs_This_stuffs_ �U  ��Y�U  ��Y�U   �Y�U  ��Y�U  A�#q�  �� /       Some_stuffs xY�U  �xY�U  �|YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0�Y�U  7E�q�  " /      Meeting     @�\�U  ��\�U  @�\Some_stuffs_Some_stuffs_ �U  ��\�U  ��\�U   �\�U  ��\�U  +�q�  � /       Meeting     Pu[�U  �u[�U  Pv[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�[�U  �q�  _ /       Meeting �U  ��\�U   �\�U  ��\Some_stuffs_Some_stuffs_ �U  �\�U  ��\�U  �\�U  ��\�U  �u�q�  A /       Appointment ��X�U  @�X�U   Yjustforfun_justforfun_ Y�U  PY�U  Y�U   	Y�U  �	Y�U  ���q�   /       Some_stuffs �O_�U  `P_�U  �P_Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   U_�U  ��>r�  (? /      Some_stuffs �x\�U  @y\�U  �y\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �}\�U  )�Jr�  IB /       Meeting �U  �^�U  �^�U  `^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �^�U  ���r�  Qe /      Some_stuffs @SZ�U   TZ�U  �TZSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  �YZ�U  A�hs�  h� /       Workout �U  �[�U  е[�U  P�[Some_stuffs_Some_stuffs_ �U  P�[�U  �[�U  й[�U  ��[�U  *�is�  �� /       Workout �U  ��[�U  P�[�U  �[justforfun_justforfun_ [�U  ��[�U  `�[�U  �\�U  P\�U  {Iks�  � /       Meeting     pH[�U  0I[�U  �I[Some_stuffs_Some_stuffs_ �U  c[�U  �c[�U  N[�U  �N[�U  $�os�  8� /      Meeting     ppZ�U  0qZ�U  p}ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0vZ�U  �t�  #� /      Workout     07[�U  �7[�U  �L[justforfun_justforfun_ _ �U  0:[�U  �:[�U  p;[�U  �;[�U  Iћ��  �( /       Meeting     �0Z�U  p1Z�U  02Zjustforfun_justforfun_ Z�U  �4Z�U  0?Z�U  7Z�U  �7Z�U  �����  Z�( /      Meeting �U  �2[�U  03[�U  �3[This_stuffs_This_stuffs_ �U  �5[�U  p6[�U  07[�U  �7[�U  �ݤ��  n�( /       Birthday    �[�U  ��[�U  ��[This_stuffs_This_stuffs_ �U  �\�U  P\�U    \�U  � \�U  e����  @%) /      Workout     `�\�U   �\�U  ��\Some_stuffs_Some_stuffs_ �U  0�\�U  ��\�U  p�\�U  ��\�U  x�Ƞ�  )) /       Appointment   Z�U  � Z�U  �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Z�U  %[��  �N) /      Workout     �w\�U   x\�U  �x\Some_stuffs_Some_stuffs_ �U   {\�U  �{\�U   |\�U  �|\�U  rp��  T) /       Birthday U  `\�U   \�U  �\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   	\�U  T��  �r) /      Meeting     �Y�U  `Y�U  �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �&Y�U  ����  �t) /       Workout �U   Z�U  �Z�U  �ZSome_stuffs_Some_stuffs_ �U  �Z�U  �Z�U  �Z�U  pZ�U  �#���  ,�) /       Workout     [�U  �[�U  P[Some_stuffs_Some_stuffs_ �U  [�U  �[�U  �[�U  P[�U  T	���  ��) /      Birthday U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  ���  ��) /       Some_stuffs 0�X�U  ��X�U  ��Xjustforfun_justforfun_ _ his_stuffs_This_stuffs_ �U  ��X�U  ���  ��) /       Workout     .\�U  �.\�U  �/\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �3\�U  
�,��  ��) /       Some_stuffs pe\�U  �e\�U  pf\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �j\�U  |B4��  ��) /      Birthday    ��[�U  P�[�U  �[Some_stuffs_Some_stuffs_ �U  г[�U  ��[�U  �[�U  е[�U  C�6��  h�) /       Birthday    �O\�U  PP\�U  �P\This_stuffs_This_stuffs_ �U  S\�U  �S\�U  PT\�U  �T\�U  h����  �) /       Appointment �<Z�U  P=Z�U  >Zjustforfun_justforfun_ Z�U  PAZ�U  �AZ�U  �BZ�U  PCZ�U  1�H��  ~* /       Appointment @�]�U  ��]�U  @�]This_stuffs_This_stuffs_ �U  @�]�U   �]�U  ��]�U  @�]�U  *d��  �* /       Meeting     �!Z�U  @"Z�U   #ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P(Z�U  se��  �* /       Workout     @SZ�U   TZ�U  �TZjustforfun_justforfun_ Z�U  �WZ�U  @XZ�U   YZ�U  �YZ�U    k��  T* /       Birthday fs ��\�U  `�\�U   �\justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  `�\�U  �d��  �6* /       Meeting                        Some_stuffs_Some_stuffs_                                     ���  �6* /       Workout     @�\�U  ��\�U  @�\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��\�U  `���  �6* /       Some_stuffs EY�U  �EY�U  �HYThis_stuffs_This_stuffs_ �U  �PY�U  @QY�U  0TY�U   VY�U  �b��  e7* /       Birthday    ppZ�U  0qZ�U  p}ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0vZ�U  ����  `;* /       Meeting     Pv[�U  w[�U  �w[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0|[�U  �����  �;* /       Meeting     pd\�U  �d\�U  pe\justforfun_justforfun_ \�U  �g\�U  0h\�U  �h\�U  �i\�U  !T���  =* /      Appointment �v\�U   w\�U  �w\justforfun_justforfun_ \�U  �y\�U  �z\�U   {\�U  �{\�U  9ꖥ�  d* /       Some_stuffs p?[�U  �?[�U  p@[justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  �D[�U  �x���  yd* /       Appointment  Z�U  �Z�U  �ZSome_stuffs_Some_stuffs_ �U  �Z�U  �Z�U  �Z�U  pZ�U  ����  ��* /       Workout     ��X�U  ��X�U  0�XSome_stuffs_Some_stuffs_ �U   �X�U  ��X�U  ��X�U  @�X�U  �U��  p�* /       Appointment ��[�U  0�[�U  �[Some_stuffs_Some_stuffs_ �U  p�[�U  0�[�U  �[�U  p�[�U  h�(��  q�* /       Meeting �U   Z�U  �Z�U  �Zjustforfun_justforfun_ Z�U  �Z�U  �Z�U  �Z�U  pZ�U  a����  ��* /       Some_stuffs �[�U  е[�U  P�[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��[�U  N����  ��* /      Workout     0�Z�U  ��Z�U  p�ZThis_stuffs_This_stuffs_ �U  0�Z�U  ��Z�U  p�Z�U  0�Z�U  �C���  ��* /       Meeting �U  ��[�U  p�[�U  0�[This_stuffs_This_stuffs_ �U  0�[�U  ��[�U  0�[�U  ��[�U  a�P��  <�* /       Meeting     �~Z�U  0Z�U  �ZThis_stuffs_This_stuffs_ �U  ��Z�U  ��Z�U  p�Z�U  0�Z�U  �WU��  \�* /      Birthday    @i[�U  �i[�U  @j[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �n[�U  a����  ��* /       Workout     ��Z�U  `�Z�U   �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ` [�U  � ���  �+ /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �&w��  � + /       Some_stuffs `�Z�U   �Z�U  оZjustforfun_justforfun_ Z�U  ��Z�U  p�Z�U  0�Z�U  ��Z�U  �ބ��  $+ /      Workout      �Y�U  ��Y�U  ��YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Z�U  ����  $+ /       Workout     P�Y�U  �Y�U  ��YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  ���  �J+ /      Appointment �Z�U  pZ�U  0	ZSome_stuffs_Some_stuffs_ �U  �Z�U  �Z�U  �Z�U  @Z�U  d����   n+ /      Meeting     0)[�U  �)[�U  �*[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p/[�U  qs���  �q+ /       Appointment P�[�U  �[�U  й[Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  ��[�U  �@��  ��+ /       Meeting  fs �%Y�U  �&Y�U  )YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �5Y�U  B�H��  ȗ+ /       Some_stuffs �a[�U  0b[�U  Pz[justforfun_justforfun_ [�U  �e[�U   f[�U  �f[�U  @g[�U  ��P��  ڙ+ /       Some_stuffs 0TY�U   VY�U  @YYThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `fY�U  �xS��  }�+ /      Birthday                       justforfun_justforfun_                                       5pU��  ��+ /       Appointment �zZ�U  �{Z�U  p|ZSome_stuffs_Some_stuffs_ �U  �Z�U  ��Z�U  p�Z�U  0�Z�U  4:^��  >�+ /       Some_stuffs @�\�U   �\�U  ��\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��\�U  n�^��  Q�+ /       Some_stuffs �eY�U  `fY�U  �iYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �xY�U  �۪�  0�+ /       Workout      �Y�U  ��Y�U  ��Yjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ��Y�U  ����  E�+ /      Workout     �eY�U  `fY�U  �iYSome_stuffs_Some_stuffs_ �U  �sY�U  `tY�U  xY�U  �xY�U  ��|��  ��+ /      Birthday    0:[�U  �:[�U  p;[This_stuffs_This_stuffs_ �U  �=[�U  �>[�U  p?[�U  �?[�U  �ď��  v�+ /       Workout �U  ��X�U  @�X�U   YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �	Y�U  �_��  V
, /       Meeting     ��Z�U  ��Z�U  @�ZThis_stuffs_This_stuffs_ �U  `�Z�U   �Z�U  ��Z�U  `�Z�U  �u	��  �
, /      Workout ffs   Z�U  � Z�U  �!ZSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  �&Z�U  �)��  �, /       Workout     ��[�U  ��[�U  @�[This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ��[�U  �栬�  b1, /       Appointment �^�U  ��^�U  �^Some_stuffs_Some_stuffs_ �U  ��^�U   �^�U  ��^�U   �^�U  1ѡ��  �1, /       Meeting     �/[�U  p0[�U  01[This_stuffs_This_stuffs_ �U  �3[�U  p4[�U  �4[�U  p5[�U  ���  7, /      Some_stuffs �[�U  0�[�U  ��[justforfun_justforfun_ _ �U  p�[�U  0�[�U  ��[�U  0�[�U   :��  �X, /       Some_stuffs `�Z�U   �Z�U  ��Zjustforfun_justforfun_ Z�U  ��Z�U  p�Z�U  0�Z�U  ��Z�U  ��B��  �Z, /      Meeting ent &Z�U  �&Z�U  �'Zjustforfun_justforfun_ _This_stuffs_This_stuffs_ �U  �,Z�U  CD��  ([, /       Some_stuffs �~Z�U  0Z�U  �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0�Z�U  2iY��  �`, /       Appointment ��Z�U  p�Z�U  0�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  ���  )�, /      Birthday    @i[�U  �i[�U  @j[This_stuffs_This_stuffs_ �U  �l[�U   m[�U  �m[�U  �n[�U  �o��  ��, /       Birthday    0_[�U  �_[�U  p`[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �d[�U   .s��  ��, /       Meeting     �zZ�U  �{Z�U  p|ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0�Z�U  �i��  ��, /       Some_stuffs ��Y�U  �Y�U  ��YThis_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  @�Y�U  �
��  ��, /      Some_stuffs ��Z�U  `�Z�U   �Zjustforfun_justforfun_ Z�U  ��Z�U  ��Z�U  0�Z�U  ��Z�U  ��G��  � - /      Meeting     0_[�U  �_[�U  p`[Some_stuffs_Some_stuffs_ �U  Pz[�U  �z[�U  @d[�U  �d[�U  P4H��  � - /       Birthday    ��Y�U  p�Y�U  ��YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Y�U  �}L��  �!- /       Workout     p@[�U  �@[�U  �A[This_stuffs_This_stuffs_ �U  0D[�U  �D[�U  �E[�U  0F[�U  �̰�  �B- /       Some_stuffs �%Y�U  �&Y�U  )YSome_stuffs_Some_stuffs_ �U  �1Y�U  �2Y�U  5Y�U  �5Y�U  ��հ�  E- /      Appointment @�[�U   �[�U   �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �[�U  ��w��  }n- /      Birthday    ��Z�U  0�Z�U  �Zjustforfun_justforfun_ Z�U  ��Z�U  0�Z�U  �Z�U  ��Z�U  z�!��  �8 /       Birthday fs �C]�U  D]�U  �D]justforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U  0H]�U  ;z5��  8 /       Birthday    @�]�U  ��]�U  `�]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p�]�U  �18��  �8 /       Workout     @ \�U  � \�U  @!\This_stuffs_This_stuffs_ �U  �#\�U  P$\�U  �$\�U  P%\�U  ��9��  :8 /      Workout     `[�U   [�U  �[This_stuffs_This_stuffs_ �U  `	[�U   
[�U  �
[�U   [�U  �Z���  �?8 /      Meeting     �+\�U  P,\�U  �,\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �1\�U  )#���  	@8 /       Some_stuffs ��]�U  `�]�U  ��]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��]�U  a�_��  |j8 /       Birthday U  PG_�U  �G_�U  PH_This_stuffs_This_stuffs_ �U  �J_�U   K_�U  �K_�U   L_�U  P>b��  k8 /       Meeting     ��Y�U  `�Y�U   �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  Z<���  ��8 /       Workout     p
Z�U  0Z�U  �Zjustforfun_justforfun_ Z�U  PZ�U  Z�U  �Z�U  �Z�U  p����  ��8 /       Appointment 7Z�U  �7Z�U  P8ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P=Z�U  n���  C�8 /      Some_stuffs p�[�U  0�[�U  ��[Some_stuffs_Some_stuffs_ �U  0�[�U  ��[�U  ��[�U  p�[�U  ���  ��8 /       Some_stuffs p{[�U  0|[�U  �|[justforfun_justforfun_ [�U  �[�U  0�[�U  ��[�U  p�[�U  5���  ¶8 /      Workout �U  @�[�U  ��[�U  @�[justforfun_justforfun_ [�U  ��[�U  @�[�U   �[�U  ��[�U  �I���  k�8 /       Birthday    P�Y�U  �Y�U  ��Yjustforfun_justforfun_ Y�U   �Y�U  ��Y�U  ��Y�U  ��Y�U  �)���  o�8 /       Meeting      Z�U  �Z�U  �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  pZ�U  [���  '�8 /       Workout     ��]�U   �]�U  ��]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P�]�U  ]a"��  ��8 /      Birthday U  P�[�U  п[�U  ��[Some_stuffs_Some_stuffs_ �U  ��[�U  P�[�U  �[�U  ��[�U  b9��  ��8 /       Meeting ffs  	Y�U  �	Y�U  �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `Y�U  X�9��  ��8 /       Appointment �Z�U  ��Z�U  @�Zjustforfun_justforfun_ Z�U  ��Z�U  ��Z�U  p�Z�U  ��Z�U  ܺV��  �,9 /      Some_stuffs �Q[�U  pR[�U  0S[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �W[�U  ��k��  #29 /       Some_stuffs ��Y�U  ��Y�U  �Yjustforfun_justforfun_ Y�U  `�Y�U   �Y�U  ��Y�U  `�Y�U  ����  /R9 /       Appointment ��Y�U  `�Y�U   �YSome_stuffs_Some_stuffs_ �U  p�Y�U  0�Y�U  ��Y�U  ��Y�U  �����  �W9 /      Meeting �U  p3Z�U  04Z�U  �4ZThis_stuffs_This_stuffs_ �U  P8Z�U  9Z�U  �9Z�U  P:Z�U  z����  �W9 /       Birthday    `E^�U  F^�U  �F^This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  J^�U  Ǆ��  z9 /      Birthday    0�[�U  �[�U  p�[Some_stuffs_Some_stuffs_ �U  0�[�U  ��[�U  0�[�U  ��[�U  P����  �}9 /       Birthday    P�\�U  Н\�U  ��\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��\�U  T� ��  ��9 /      Some_stuffs  �Y�U  �Y�U  0�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Y�U  �y"��  m�9 /       Birthday    p�]�U  �]�U  ��]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �]�U  `���  �9 /       Meeting      �\�U  ��\�U   �\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �\�U  �JV��  :�9 /       Workout     EY�U  �EY�U  �HYThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   VY�U  �sb��  W�9 /       Workout     0�Z�U  ��Z�U  p�ZSome_stuffs_Some_stuffs_ �U  ��Z�U  ��Z�U  0�Z�U  � [�U  4����  �: /      Birthday                       justforfun_justforfun_                                       �[���  �: /       Meeting     ��Y�U  ��Y�U  p�YSome_stuffs_Some_stuffs_ �U  ��Y�U  @�Y�U   �Y�U  ��Y�U  4����  b?: /      Appointment �QZ�U  �RZ�U  �HZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �MZ�U  �r���  eA: /       Birthday    ��Y�U  `�Y�U   �YThis_stuffs_This_stuffs_ �U  p�Y�U  0�Y�U  ��Y�U  ��Y�U  �w��  �c: /      Workout                        This_stuffs_This_stuffs_                                     ��$��  �g: /       Some_stuffs  �]�U  ��]�U   �]justforfun_justforfun_ _ �U   �]�U  ��]�U   �]�U  ��]�U  �&��  �g: /       Workout     ��Y�U  ��Y�U   �YSome_stuffs_Some_stuffs_ �U  ��Y�U  ��Y�U   �Y�U  ��Y�U  +�*��  )i: /       Workout     �J^�U  PK^�U  �K^Some_stuffs_Some_stuffs_ �U  N^�U  �N^�U  O^�U  �O^�U  @����  h�: /       Workout     �[�U  �[�U  [Some_stuffs_Some_stuffs_ �U  �[�U  �[�U  P[�U  [�U  �����  ��: /      Meeting     ��^�U  `�^�U  ��^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��^�U  fF��  ı: /      Birthday    �zZ�U  �{Z�U  p|ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0�Z�U  P���  r�: /       Appointment `\�U   \�U  �\Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   	\�U  �kw��  ��: /      Workout     �W^�U  PX^�U  �X^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �\^�U  PȌ��  R; /       Workout �U  p^�U  �^�U  p^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0"^�U  
Q
��  u%; /       Workout     �rZ�U  psZ�U  0tZThis_stuffs_This_stuffs_ �U  �vZ�U  pwZ�U  0xZ�U  �xZ�U  �>��  �*; /       Birthday    ��Z�U  `�Z�U   �Zjustforfun_justforfun_ Z�U  `�Z�U   �Z�U  ��Z�U  ��Z�U  55,��  ".; /      Workout     �%Y�U  �&Y�U  )YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �5Y�U  ���  �S; /      Meeting     И]�U  P�]�U  Й]This_stuffs_This_stuffs_ �U  Л]�U  ��]�U   �]�U  ��]�U  @����  hT; /       Workout     �Z�U  �Z�U  �ZThis_stuffs_This_stuffs_ �U  p
Z�U  0Z�U  �Z�U  �Z�U  D+C��  �u; /      Some_stuffs                    justforfun_justforfun_                                       acD��  �u; /       Workout     5Y�U  �5Y�U  P8YThis_stuffs_This_stuffs_ �U  @?Y�U  AY�U  EY�U  �EY�U  �I��  w; /       Workout     �QZ�U  �RZ�U  �HZSome_stuffs_Some_stuffs_ �U  �KZ�U  pLZ�U  0MZ�U  �MZ�U  �*R��  cy; /       Meeting ent pP[�U  0Q[�U  �Q[justforfun_justforfun_ _ �U  pT[�U  �T[�U  �U[�U  0V[�U  �c���  ��; /       Birthday    �k]�U  @l]�U  �l]This_stuffs_This_stuffs_ �U   o]�U  �o]�U  @p]�U  �p]�U  t���  Y�; /      Workout     @�Z�U  ��Z�U  �ZThis_stuffs_This_stuffs_ �U  p�Z�U  ��Z�U  ��Z�U  p�Z�U  )j���  i�; /       Workout ffs �Q]�U  pR]�U  �$]justforfun_justforfun_ _ �U  �&]�U  �']�U  @(]�U  �(]�U  ��m��  �; /      Appointment Pu[�U  �u[�U  Pv[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�[�U  �v��  �; /       Some_stuffs  j\�U  �j\�U  @k\justforfun_justforfun_ \�U  �m\�U   n\�U  �n\�U  @o\�U  �|��  ��; /       Appointment �zZ�U  �{Z�U  p|ZThis_stuffs_This_stuffs_ �U  �Z�U  ��Z�U  p�Z�U  0�Z�U  ����  k�; /       Workout     7Z�U  �7Z�U  P8Zjustforfun_justforfun_ Z�U  ;Z�U  �;Z�U  �<Z�U  P=Z�U  �,��  ��; /       Birthday nt s[�U  �s[�U  t[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Px[�U  �"��  %�; /       Birthday U  �|]�U   }]�U  �}]This_stuffs_This_stuffs_ �U   �]�U  ��]�U  0�]�U  ��]�U  ��(��  ��; /       Meeting      �Z�U  ��Z�U  0�Zjustforfun_justforfun_ _ �U  0�Z�U  ��Z�U  p�Z�U  ��Z�U  lf���  �< /      Appointment ppZ�U  0qZ�U  p}ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0vZ�U  ᧴��  �< /       Workout ffs `�Y�U   �Y�U  ��YThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  0�Y�U  �`x��  P�< /      Appointment �%Y�U  �&Y�U  )YThis_stuffs_This_stuffs_ �U  �1Y�U  �2Y�U  5Y�U  �5Y�U  ���  �[G /       Some_stuffs �[�U  л[�U  P�[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �[�U  ����  X^G /       Birthday    �[�U  ��[�U  ��[justforfun_justforfun_ [�U  �[�U  ��[�U  ��[�U  �[�U  .���  �`G /      Meeting     P8Z�U  9Z�U  �9ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pHZ�U  e�S�  ��G /       Meeting     ��Z�U   �Z�U   �ZThis_stuffs_This_stuffs_ �U  `�Z�U   �Z�U  ��Z�U  `�Z�U  �T�  .�G /      Birthday    �f[�U  @g[�U   h[This_stuffs_This_stuffs_ �U  @j[�U  �j[�U  @k[�U  �k[�U  4'Y�  ^�G /       Birthday fs 0�Z�U  ��Z�U  p�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Z�U  Y�\�  G�G /       Meeting     �jZ�U  pkZ�U  0lZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0qZ�U  ;�g�  �G /       Birthday    ��[�U  `�[�U  �\This_stuffs_This_stuffs_ �U  `\�U  �\�U  `\�U  �\�U  �m�  ��G /       Birthday    ppZ�U  0qZ�U  p}Zjustforfun_justforfun_ Z�U  0tZ�U  �tZ�U  puZ�U  0vZ�U  0��  ~�G /       Birthday    �J\�U  PK\�U  L\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  PP\�U  pݢ�  ��G /       Birthday    �HY�U  �IY�U  �LYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ZY�U  ���  ��G /      Appointment ��[�U  ��[�U  @�[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��[�U  y#�  ��G /       Workout      �[�U  ��[�U  ��[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �[�U  �:1�  8�G /       Meeting     ��[�U  ��[�U  �[justforfun_justforfun_ [�U  ��[�U  P�[�U  �[�U  ��[�U  L���  �H /      Appointment 0TY�U   VY�U  @YYThis_stuffs_This_stuffs_ �U  paY�U  0bY�U  �eY�U  `fY�U  �=��  �!H /       Meeting     @A\�U   B\�U  �B\Some_stuffs_Some_stuffs_ �U  0E\�U  �E\�U  PF\�U  G\�U  �V]�  IH /       Some_stuffs 0�[�U  ��[�U  ��[justforfun_justforfun_ [�U  ��[�U  p�[�U  0�[�U  ��[�U  �ic�  �JH /      Some_stuffs @�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_ �U  ��Z�U  `�Z�U   �Z�U  ��Z�U  pg��  rH /       Appointment �h\�U  �i\�U   j\This_stuffs_This_stuffs_ �U  @l\�U  �l\�U  �m\�U   n\�U  �҈�  ��H /       Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             Ka��  �H /       Appointment ��\�U  ��\�U  @�\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �\�U  ]���  K�H /      Meeting       Z�U  � Z�U  �!ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �&Z�U  ���  O�H /       Workout     �\�U  @>\�U  \Some_stuffs_Some_stuffs_ �U  @!\�U  �!\�U  p"\�U  �"\�U  ��"�  #�H /       Some_stuffs PS^�U  �S^�U  �T^This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  PX^�U  �\'�  M�H /       Some_stuffs оZ�U  P�Z�U  0�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Z�U  ݁*�  �H /      Some_stuffs �'Z�U  P(Z�U  )ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P6Z�U  ,p6�  )�H /       Workout     �^�U  `^�U  �^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �^�U  ;9�  ��H /       Meeting     �\�U  p\�U  0\Some_stuffs_Some_stuffs_ �U  p\�U  �\�U  �\�U  p\�U  +��  ��H /      Birthday    @�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  A���  h�H /       Appointment �]�U  �]�U  0]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0]�U  �1��  D�H /       Birthday    �[�U  е[�U  P�[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��[�U  "�J�  �I /       Birthday    �yZ�U  0zZ�U  �zZjustforfun_justforfun_ Z�U  �~Z�U  0Z�U  �Z�U  ��Z�U  lP�  Y
I /      Birthday                       Some_stuffs_Some_stuffs_                                     �0R�  �
I /       Meeting     @ \�U  � \�U  @!\Some_stuffs_Some_stuffs_ �U  �#\�U  P$\�U  �$\�U  P%\�U  �i^�  �I /       Meeting     `�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_ �U  ��Z�U  ��Z�U  @�Z�U   �Z�U  �^��  �4I /      Workout     p�Z�U  0�Z�U  ��ZThis_stuffs_This_stuffs_ �U  0�Z�U  �Z�U  ��Z�U  0�Z�U  (r}�  iWI /       Meeting      �Z�U  ��Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �Z�U  uj�  �WI /      Meeting     )Z�U  �)Z�U  P*ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �.Z�U  l��  1~I /       Appointment 0)[�U  �)[�U  �*[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p/[�U  b�#�  ��I /       Appointment 0MZ�U  �MZ�U  pNZSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   TZ�U  �<*�  ��I /       Birthday U  @SZ�U   TZ�U  �TZThis_stuffs_This_stuffs_ �U  �WZ�U  @XZ�U   YZ�U  �YZ�U  �+�  ڃI /       Meeting �U  �F]�U  0G]�U  �G]justforfun_justforfun_ ]�U  �I]�U  �J]�U  K]�U  �K]�U  -&3�  �I /      Some_stuffs  �Y�U  �Y�U  0�Yjustforfun_justforfun_ Y�U  ��Y�U  ��Y�U  P�Y�U  �Y�U  ~��  ?�I /       Appointment �<Z�U  P=Z�U  >Zjustforfun_justforfun_ Z�U  PAZ�U  �AZ�U  �BZ�U  PCZ�U  �o��  שI /       Appointment ppZ�U  0qZ�U  p}Zjustforfun_justforfun_ Z�U  0tZ�U  �tZ�U  puZ�U  0vZ�U  N���  A�I /      Workout     @k[�U  �k[�U  �l[Some_stuffs_Some_stuffs_ �U   o[�U  �o[�U  @p[�U   q[�U  ��K �  ��I /       Some_stuffs @k[�U  �k[�U  �l[Some_stuffs_Some_stuffs_ �U   o[�U  �o[�U  @p[�U   q[�U  �zQ �  :�I /      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��Y �  Y�I /       Some_stuffs ppZ�U  0qZ�U  p}ZThis_stuffs_This_stuffs_ �U  0tZ�U  �tZ�U  puZ�U  0vZ�U  ��� �  =�I /      Birthday    0TY�U   VY�U  @YYjustforfun_justforfun_ Y�U  paY�U  0bY�U  �eY�U  `fY�U  I�w!�  �J /       Workout     p3Z�U  04Z�U  �4ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P:Z�U  h݈!�  �J /       Appointment  �Y�U  ��Y�U  ��YSome_stuffs_Some_stuffs_ �U  �Z�U  `Z�U   Z�U  �Z�U  �k�!�  �J /      Appointment 0]�U  �]�U  p	]Some_stuffs_Some_stuffs_ �U  �]�U  �]�U  0]�U  �]�U  ��"�  �@J /       Appointment �.]�U  �/]�U  0]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �3]�U  �!"�  $FJ /      Some_stuffs xY�U  �xY�U  �|YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0�Y�U  �""�  -FJ /       Workout     p�Y�U  0�Y�U  0�YThis_stuffs_This_stuffs_ �U   �Y�U  ��Y�U  ��Y�U  p�Y�U  �"�  �gJ /       Meeting ent �]Z�U  `^Z�U   _ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `dZ�U  j��"�  �oJ /       Workout     �?Z�U  �@Z�U  PAZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  PFZ�U  9;�"�  �pJ /       Birthday    0D[�U  �D[�U  �E[This_stuffs_This_stuffs_ �U  pH[�U  0I[�U  �I[�U  pJ[�U  ��A#�  ׏J /       Some_stuffs �%]�U  p&]�U  �&]justforfun_justforfun_ ]�U  p)]�U  �)]�U  p*]�U   +]�U  J>K#�  =�J /       Meeting     �WZ�U  @XZ�U   YZSome_stuffs_Some_stuffs_ �U   \Z�U  pgZ�U  �]Z�U  `^Z�U  Xd`#�  ��J /       Meeting     02Z�U  �2Z�U  p3ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  9Z�U  �b�#�  <�J /      Appointment  Z�U  �Z�U  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pZ�U  �$�  �J /      Appointment �Z�U  @Z�U  PZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  PZ�U  �%�  $K /       Some_stuffs ��Z�U  ��Z�U  @�ZSome_stuffs_Some_stuffs_ �U   �Z�U  ��Z�U  ��Z�U   �Z�U  �P�%�  �-K /      Appointment ��[�U  P�[�U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P�[�U  �c�%�  �-K /       Appointment 0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  ��X�U  ��%�  �1K /       Appointment �9]�U  �:]�U   ;]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `?]�U  +O>&�  �SK /       Appointment �\�U  p\�U  0\Some_stuffs_Some_stuffs_ �U  �\�U  p\�U  0\�U  �\�U  H�>&�  �SK /       Workout �U    Z�U  � Z�U  �!ZSome_stuffs_Some_stuffs_ �U  �$Z�U  p-Z�U  &Z�U  �&Z�U  ��H&�  CVK /       Appointment �;Y�U  `<Y�U  @?YSome_stuffs_Some_stuffs_ �U  �HY�U  �IY�U  �LY�U  `MY�U  e�R&�  �XK /      Meeting      �Y�U  ��Y�U  ��Yjustforfun_justforfun_ Y�U  P�Y�U  �Y�U  ��Y�U  ��Y�U  ҅�&�  �zK /       Workout ent ��Z�U  ��Z�U  @�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  y��&�  ~K /       Some_stuffs �[^�U  �\^�U  0]^Some_stuffs_Some_stuffs_ �U  `_^�U  ��^�U  ``^�U  a^�U  ��&�  C�K /       Workout     оZ�U  P�Z�U  0�ZSome_stuffs_Some_stuffs_ �U  0�Z�U  ��Z�U  0�Z�U  �Z�U  0�o'�  ��K /       Some_stuffs   Z�U  � Z�U  �!ZThis_stuffs_This_stuffs_ �U  �$Z�U  p-Z�U  &Z�U  �&Z�U  ��s'�  ͢K /       Birthday      \�U  � \�U  `\Some_stuffs_Some_stuffs_ �U  `\�U   \�U  �\�U   \�U  �}'�  N�K /      Meeting     )Z�U  �)Z�U  P*ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �.Z�U  cf'�  ��K /       Meeting ent �y\�U  �z\�U   {\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �~\�U  N(�  ?�K /       Appointment P�Y�U  �Y�U  ��YSome_stuffs_Some_stuffs_ �U   �Y�U  ��Y�U  ��Y�U  ��Y�U  �h(�  ��K /      Meeting     ��X�U  ��X�U  0�XSome_stuffs_Some_stuffs_ �U   �X�U  ��X�U  ��X�U  @�X�U  (�  x�K /       Workout     �4Z�U  0?Z�U  7ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �;Z�U  |ۦ(�  _�K /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �*TR�  ��V /       Workout     .\�U  �.\�U  �/\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �3\�U  ЛrR�  ��V /       Some_stuffs p%[�U  0&[�U  �&[This_stuffs_This_stuffs_ �U  0)[�U  �)[�U  �*[�U  p+[�U   ��R�  ��V /       Workout     02Z�U  �2Z�U  p3ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  9Z�U  ��R�  /�V /       Some_stuffs P�[�U  з[�U  P�[Some_stuffs_Some_stuffs_ �U  �[�U  л[�U  P�[�U  �[�U  �ˑS�  �V /      Birthday     �Y�U  ��Y�U  ��YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  9�S�  ��V /       Birthday nt  �Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  p�Z�U   g�T�  �9W /       Some_stuffs �P\�U  PQ\�U  �Q\Some_stuffs_Some_stuffs_ �U  PT\�U  �T\�U  PU\�U  �U\�U  i�T�  J=W /       Appointment �%Y�U  �&Y�U  )YThis_stuffs_This_stuffs_ �U  �1Y�U  �2Y�U  5Y�U  �5Y�U  �pU�  xhW /       Workout     �Z�U  pZ�U  0	ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @Z�U  ��U�  όW /       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �V�  ^�W /      Workout     @�[�U  ��[�U  ��[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �[�U  (��V�  ɯW /       Workout �U  0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��X�U  :��V�  S�W /       Appointment �Z�U  `�Z�U  �Zjustforfun_justforfun_ Z�U  `�Z�U   �Z�U  оZ�U  P�Z�U  �ʐV�  a�W /       Meeting     �Z�U  �%Z�U  �ZThis_stuffs_This_stuffs_ �U  �!Z�U  @"Z�U   #Z�U  �#Z�U  cE W�  �W /       Workout     0�\�U  ��\�U  p�\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P�\�U  �b,W�  6�W /       Meeting     ��[�U  `�[�U  �\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �\�U  ��,W�  Z�W /      Birthday      ]�U  � ]�U  0!]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pR]�U  ��2W�  ��W /       Some_stuffs `�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �Z�U  Y�2W�  ��W /       Appointment ��[�U  0�[�U  �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�[�U  �=<W�  E�W /       Some_stuffs ��[�U  @�[�U   �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��[�U  ��W�  �W /       Birthday     (^�U  �(^�U   )^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �,^�U  `[�W�  � X /       Appointment 0�X�U  ��X�U  ��Xjustforfun_justforfun_ X�U  ��X�U  ��X�U  ��X�U  ��X�U  R��X�  rJX /       Some_stuffs �m\�U   n\�U  �n\justforfun_justforfun_ _ his_stuffs_This_stuffs_ �U  @s\�U  ���X�  �LX /       Workout     ��Z�U  `�Z�U   �Zjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ��Z�U   ?�X�  `MX /       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             յ�X�  �NX /      Workout ent ��X�U  @�X�U   Yjustforfun_justforfun_ Y�U  PY�U  Y�U   	Y�U  �	Y�U  Ln�X�  =PX /       Some_stuffs @�\�U  ��\�U  @�\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��\�U  ��Y�  5vX /       Workout     `�Z�U   �Z�U  �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �Z�U  ��Z�  �X /       Some_stuffs                    Some_stuffs_Some_stuffs_                                     �Z�  Y�X /      Appointment p�Z�U  0�Z�U   �ZThis_stuffs_This_stuffs_ �U  ��Z�U  p�Z�U  0�Z�U  ��Z�U  C˻Z�  ��X /       Some_stuffs ��Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_ �U  ��Z�U  @�Z�U   �Z�U  ��Z�U  �.�Z�  ��X /       Meeting �U   _Z�U  �_Z�U  �`ZSome_stuffs_Some_stuffs_ �U  �cZ�U  `dZ�U   eZ�U  �eZ�U  9[�Z�  ��X /       Birthday    p;[�U  �;[�U  �<[Some_stuffs_Some_stuffs_ �U  p?[�U  �?[�U  p@[�U  �@[�U  v�Z�  ��X /      Workout     0�[�U  Ь[�U  0�[This_stuffs_This_stuffs_ �U  �[�U  ��[�U  0�[�U  �[�U  (N[�   �X /       Workout     ��Z�U  ��Z�U  @�ZThis_stuffs_This_stuffs_ �U  @�Z�U   �Z�U  ��Z�U  ��Z�U  ��X[�  ��X /       Meeting      	Y�U  �	Y�U  �YThis_stuffs_This_stuffs_ �U  �Y�U  `Y�U  �Y�U  `Y�U  �X`[�  ��X /      Workout     �Z�U   Z�U  �ZThis_stuffs_This_stuffs_ �U  �Z�U  pZ�U  0	Z�U  �	Z�U  ��[�  LY /       Workout     ��\�U   �\�U  ��\justforfun_justforfun_ \�U  P�\�U  Щ\�U  p�\�U  0�\�U  t��[�  �Y /      Birthday U  �QZ�U  �RZ�U  �HZjustforfun_justforfun_ Z�U  �KZ�U  pLZ�U  0MZ�U  �MZ�U  �!�\�  �7Y /       Appointment EY�U  �EY�U  �HYThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   VY�U  ܷ�\�  �<Y /      Appointment xY�U  �xY�U  �|YSome_stuffs_Some_stuffs_ �U  ��Y�U  ��Y�U  p�Y�U  0�Y�U  �Z(]�  ebY /      Meeting �U  ��Z�U  p�Z�U  0�ZSome_stuffs_Some_stuffs_ �U  p�Z�U  0�Z�U  ��Z�U  0�Z�U  �,�]�  $�Y /       Workout     �P\�U  PQ\�U  �Q\Some_stuffs_Some_stuffs_ �U  PT\�U  �T\�U  PU\�U  �U\�U  �Ʊ]�  ��Y /      Birthday    `�Y�U   �Y�U  ��YSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  0�Y�U  @��]�  (�Y /       Birthday    ��Y�U  `�Y�U   �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  �,�]�  x�Y /       Workout     0\�U  �\�U  �\justforfun_justforfun_ \�U  �\�U  p\�U  0\�U  �\�U  ���]�  %�Y /       Birthday    И]�U  P�]�U  Й]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��]�U  ��?^�  ��Y /       Appointment �Z�U  @Z�U  PZSome_stuffs_Some_stuffs_ �U  PZ�U  �Z�U  �Z�U  PZ�U  ��@^�  ;�Y /      Some_stuffs �gZ�U  phZ�U  0iZjustforfun_justforfun_ Z�U  0lZ�U  �lZ�U  pmZ�U  0nZ�U  j
L^�  �Y /       Appointment 0�[�U  ��[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0�[�U  ��^�  2�Y /      Appointment ��Y�U  ��Y�U  �YThis_stuffs_This_stuffs_ �U  `�Y�U   �Y�U  ��Y�U  `�Y�U  �xx_�  ��Y /       Birthday    @ \�U  � \�U  @!\This_stuffs_This_stuffs_ �U  �#\�U  P$\�U  �$\�U  P%\�U  ��~_�  ��Y /       Workout     �A[�U  0B[�U  �B[Some_stuffs_Some_stuffs_ �U  �E[�U  0F[�U  �F[�U  �G[�U  N�_�  ��Y /       Some_stuffs �v]�U  �w]�U   x]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   |]�U  �m�_�  ��Y /      Meeting      _Z�U  �_Z�U  �`ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �eZ�U  Į`�  �"Z /      Birthday     h[�U  �h[�U  @i[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   m[�U  �ڦ`�  cGZ /       Appointment ��Y�U   �Y�U  ��YThis_stuffs_This_stuffs_ �U  ��Y�U  ��Y�U  �Y�U  ��Y�U  ���`�  %KZ /      Birthday fs 0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  2ظ`�  �KZ /       Workout     �Y�U  @ Y�U  �"YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0.Y�U  a5�`�  MZ /       Workout     �0Z�U  p1Z�U  02ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �7Z�U  �v�`�  �NZ /       Appointment �B[�U  pC[�U  0D[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0I[�U  ��:a�  LmZ /       Birthday     �\�U  ��\�U   �\Some_stuffs_Some_stuffs_ �U  ��\�U  p$]�U  ��\�U  ��\�U  �!Xa�  �tZ /       Appointment �L[�U  pM[�U  �8[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p=[�U  �]a�  .vZ /      Birthday    �Z�U  �Z�U  `Zjustforfun_justforfun_ Z�U  �Z�U  @Z�U    Z�U  � Z�U  ���a�  ��Z /      Workout     @t]�U  �t]�U  @u]Some_stuffs_Some_stuffs_ �U   x]�U  �x]�U   y]�U  �y]�U  H��a�  ��Z /       Birthday U  P�Y�U  �Y�U  ��YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  ��zb�  /�Z /       Workout     @k[�U  �k[�U  �l[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   q[�U  ���b�  E�Z /      Birthday    [�U  �[�U  P[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P[�U  �A�b�  k�Z /       Meeting      {\�U  �{\�U   |\This_stuffs_This_stuffs_ �U  @~\�U  �~\�U  @\�U  �\�U  �_c�  ��Z /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             1&c�  ��Z /       Workout     ��X�U  @�X�U   YSome_stuffs_Some_stuffs_ �U  PY�U  Y�U   	Y�U  �	Y�U  
J�c�  [ /       Some_stuffs 0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  ֧c�  ?[ /       Workout     p�Z�U  �Z�U  ��ZThis_stuffs_This_stuffs_ �U  @�Z�U   �Z�U  ��Z�U  ��Z�U  `òc�  [ /      Birthday U  0�[�U  ��[�U  ��[This_stuffs_This_stuffs_ �U  0�[�U  Ь[�U  0�[�U  �[�U  8еc�  �[ /       Some_stuffs p�Y�U  0�Y�U  ��Yjustforfun_justforfun_ Y�U  ��Y�U  ��Y�U   �Y�U  ��Y�U  Ҷc�  [ /       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �V�c�  7[ /       Appointment  �Y�U  ��Y�U  ��YSome_stuffs_Some_stuffs_ �U  P�Y�U  �Y�U  ��Y�U  ��Y�U  Đ��  ��e /      Appointment 0\�U  �\�U  �\justforfun_justforfun_ \�U  �\�U  0\�U  �\�U  p\�U  �����  �f /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ٶ���  7f /       Birthday    GZ�U  �GZ�U  �QZjustforfun_justforfun_ Z�U  0JZ�U  �JZ�U  �KZ�U  pLZ�U  ��!��  �-f /      Birthday fs V]�U  �V]�U  PW]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   \]�U  (A��  �5f /       Some_stuffs @�[�U   �[�U   �[justforfun_justforfun_ [�U  @�[�U  ��[�U  ��[�U  �[�U  ��B��  �5f /       Some_stuffs  �Z�U  �Z�U  `�ZThis_stuffs_This_stuffs_ �U  �Z�U  ��Z�U   �Z�U  ��Z�U  �ݹ��  rTf /      Some_stuffs  eZ�U  �eZ�U  �fZThis_stuffs_This_stuffs_ �U  0iZ�U  �iZ�U  �jZ�U  pkZ�U  i[Ώ�  �Yf /       Workout     �?Z�U  �@Z�U  PAZSome_stuffs_Some_stuffs_ �U  DZ�U  �DZ�U  �EZ�U  PFZ�U  �R��  �{f /       Appointment �Q[�U  pR[�U  0S[Some_stuffs_Some_stuffs_ �U  �U[�U  0V[�U  �V[�U  �W[�U  �Y��  3}f /      Meeting ffs �X]�U  �Y]�U  @Z]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `^]�U  ����  ȣf /      Appointment p�Y�U  0�Y�U  0�Yjustforfun_justforfun_ Y�U   �Y�U  ��Y�U  ��Y�U  p�Y�U  0n���  ��f /       Appointment                    Some_stuffs_Some_stuffs_                                     ᵆ��  l�f /       Appointment 0�[�U  ��[�U  0�[justforfun_justforfun_ [�U  p�[�U  0�[�U  ��[�U  p�[�U  `G���  \�f /       Workout �U  ppZ�U  0qZ�U  p}ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0vZ�U  �i+��  ��f /       Birthday nt �#\�U  P$\�U  �$\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �)\�U  p�2��  ��f /       Workout     ��[�U   �[�U  ��[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @�[�U  =y���  wg /      Appointment P]Y�U  ^Y�U  paYSome_stuffs_Some_stuffs_ �U  �iY�U  �jY�U  @oY�U   pY�U  hɒ�  �g /       Birthday nt p�Z�U  0�Z�U  ��ZThis_stuffs_This_stuffs_ �U  0�Z�U  �Z�U  ��Z�U  0�Z�U  �>Ӓ�  �g /       Some_stuffs @�\�U   �\�U  ��\justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ��\�U  ,�P��  �?g /      Meeting �U  @�]�U  ��]�U  @�]This_stuffs_This_stuffs_ �U  @�]�U   �]�U  ��]�U  @�]�U  QFR��  @g /       Some_stuffs 0�[�U  ��[�U  p�[justforfun_justforfun_ [�U  ��[�U  ��[�U  0�[�U  ��[�U  ;]��  �Bg /       Appointment �T]�U  �U]�U  V]justforfun_justforfun_ ]�U  �X]�U  �Y]�U  @Z]�U  �Z]�U  ���  0gg /       Meeting     �]�U  p�]�U  �]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��]�U  @Y��  Hhg /       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ]���  �kg /      Workout     `�Z�U   �Z�U  оZSome_stuffs_Some_stuffs_ �U  ��Z�U  p�Z�U  0�Z�U  ��Z�U  �q���  D�g /       Meeting �U  ��\�U  `�\�U   �\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `�\�U  �$���  x�g /       Workout �U  ��[�U  0�[�U  �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�[�U  n����  Ւg /      Appointment L]�U  �L]�U  M]This_stuffs_This_stuffs_ �U  PO]�U  �O]�U  PP]�U  �P]�U  �ѕ�  ��g /      Appointment P�Y�U  �Y�U  ��YThis_stuffs_This_stuffs_ �U   �Y�U  ��Y�U  ��Y�U  ��Y�U  ��\��  Xh /       Some_stuffs �Z�U  �%Z�U  �ZThis_stuffs_This_stuffs_ �U  �!Z�U  @"Z�U   #Z�U  �#Z�U  ��e��  �	h /      Meeting �U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  Q���  �)h /       Some_stuffs �R]�U  pS]�U  �S]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  X]�U  ����  D-h /       Appointment 0]�U  �]�U  p]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �]�U  �~���  ;/h /      Meeting     p�Z�U  0�Z�U  ��ZSome_stuffs_Some_stuffs_ �U  0�Z�U  �Z�U  ��Z�U  0�Z�U  �!z��  kPh /       Workout                        justforfun_justforfun_                                       >����  7Th /      Workout ent  
^�U  �
^�U   ^This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  �^�U  ٴ���  �Vh /       Workout     ��Y�U  ��Y�U  p�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  ���  Mwh /       Meeting                        Some_stuffs_Some_stuffs_                                     ���  Zyh /       Appointment P*\�U  +\�U  �+\Some_stuffs_Some_stuffs_ �U  .\�U  �.\�U  �/\�U  P0\�U  ����  �zh /      Birthday    ��Y�U  p�Y�U  ��YSome_stuffs_Some_stuffs_ �U  �Y�U  ��Y�U   �Y�U  �Y�U  ?Ѳ��  w�h /      Some_stuffs ��\�U  ��\�U   �\justforfun_justforfun_ \�U   �\�U  ��\�U  `�\�U   �\�U  Q����  ��h /       Birthday    ��Z�U  `�Z�U   �ZThis_stuffs_This_stuffs_ �U  `�Z�U   �Z�U  ��Z�U  ��Z�U  p
Ș�  �h /       Appointment ��Z�U  p�Z�U  0�ZSome_stuffs_Some_stuffs_ �U  ��Z�U  0�Z�U  �Z�U  ��Z�U  ro̘�  �h /       Meeting      Z�U  �Z�U  �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  pZ�U  T�A��  �h /      Birthday    ��[�U  0�[�U  �[Some_stuffs_Some_stuffs_ �U  p�[�U  0�[�U  �[�U  p�[�U  �ߙ�  v�h /       Birthday U   o[�U  �o[�U  @p[justforfun_justforfun_ [�U  s[�U  �s[�U  t[�U  �t[�U  :q��  s�h /       Birthday    @�\�U  ��\�U  p�\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Н\�U  [6��  ��h /       Appointment �^�U  ^�U  �^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `^�U  ��  `�h /       Birthday    p-[�U  �-[�U  �.[This_stuffs_This_stuffs_ �U  01[�U  �1[�U  �2[�U  03[�U  �s��  ;i /      Workout     p;[�U  �;[�U  �<[This_stuffs_This_stuffs_ �U  p?[�U  �?[�U  p@[�U  �@[�U  ��u��  �i /       Birthday    P�Y�U  �Y�U  ��YSome_stuffs_Some_stuffs_ �U   �Y�U  ��Y�U  ��Y�U  ��Y�U  ����  yi /       Appointment �=]�U   >]�U  �>]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  C]�U  ���  `?i /       Workout     �\�U  `\�U   \This_stuffs_This_stuffs_ �U  �	\�U  �
\�U   \�U  �\�U  j�#��  q@i /       Meeting      �Z�U  ��Z�U  `�Zjustforfun_justforfun_ Z�U  0�Z�U  �Z�U  ��Z�U  p�Z�U  ,*��  Bi /      Appointment p�Z�U  0�Z�U  ��ZThis_stuffs_This_stuffs_ �U  ��Z�U  ��Z�U  p�Z�U  ��Z�U  }r���  �ei /      Meeting     p�Z�U  ��Z�U  p�ZThis_stuffs_This_stuffs_ �U  0�Z�U  ��Z�U  ��Z�U  p�Z�U  Hɺ��  gi /       Appointment �Z�U  pZ�U  0	ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @Z�U  L���  �gi /       Workout     ��Z�U  ��Z�U  @�ZThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  `�Z�U  ,�>��  �i /       Some_stuffs @�[�U  ��[�U  ��[This_stuffs_This_stuffs_ �U  �[�U  ��[�U  ��[�U  P�[�U  )3C��  	�i /       Birthday nt  _Z�U  �_Z�U  �`ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �eZ�U  �W��  "�i /       Birthday nt �]�U  @]�U  �]justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  �"]�U   �\��  ��i /       Meeting     ��Y�U  ��Y�U  ��Yjustforfun_justforfun_ Y�U  ��Y�U   �Y�U  ��Y�U  ��Y�U  �7]��  ��i /      Appointment ��Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_ �U  `�Z�U   �Z�U  ��Z�U  `�Z�U  ���  �i /       Birthday nt �]�U  p�]�U   �]Some_stuffs_Some_stuffs_ �U   �]�U  ��]�U   �]�U  ��]�U  t���  j�i /      Some_stuffs ��Z�U  ��Z�U  @�ZSome_stuffs_Some_stuffs_ �U   �Z�U  ��Z�U  ��Z�U   �Z�U  9ox��  3�i /       Appointment `\�U   \�U  �\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   	\�U  �Q���  D�i /       Appointment `�\�U   �\�U  ��\justforfun_justforfun_ \�U  0�\�U  ��\�U  p�\�U  ��\�U  ތ��  n�i /      Birthday    ��Z�U  p�Z�U  0�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  M��  A�i /      Workout     p�Z�U  0�Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0�Z�U   ���  tj /       Workout     �zZ�U  �{Z�U  p|ZThis_stuffs_This_stuffs_ �U  �Z�U  ��Z�U  p�Z�U  0�Z�U  $i���  �$j /      Workout ffs �&^�U  �'^�U   (^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �+^�U  �ݾ��  �,j /       Some_stuffs �x[�U  �y[�U  ��[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �~[�U  1�B��  ~Nj /       Birthday nt �Z�U  �Z�U  �ZThis_stuffs_This_stuffs_ �U  p
Z�U  0Z�U  �Z�U  �Z�U  �E��  EOj /      Appointment ��X�U  ��X�U  0�XSome_stuffs_Some_stuffs_ �U   �X�U  ��X�U  ��X�U  @�X�U  ����  �wj /       Some_stuffs 0[[�U  �[[�U  0\[Some_stuffs_Some_stuffs_ �U  0_[�U  �_[�U  p`[�U  �`[�U  �.��  �yj /      Appointment �Y�U  `Y�U  �YSome_stuffs_Some_stuffs_ �U  �"Y�U  `#Y�U  �%Y�U  �&Y�U  �X���  �"u /      Birthday    ppZ�U  0qZ�U  p}ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0vZ�U  /�#��  �Hu /      Some_stuffs �"^�U  �_^�U  �$^This_stuffs_This_stuffs_ �U  �&^�U  �'^�U   (^�U  �(^�U  _0��  �Ku /       Appointment �2[�U  03[�U  �3[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �7[�U  :�4��  �Lu /       Appointment  �]�U  ��]�U  @�]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �]�U  Q�;��  �Nu /       Some_stuffs `�Z�U   �Z�U  ��Zjustforfun_justforfun_ Z�U  `�Z�U  ��Z�U  `�Z�U   �Z�U  �����  �ou /      Some_stuffs  �[�U  ��[�U  ��[justforfun_justforfun_ [�U  ��[�U  �[�U  ��[�U  ��[�U  ҽ��  pu /       Meeting     ��[�U  P�[�U  �[Some_stuffs_Some_stuffs_ �U  ��[�U  `�[�U   �[�U  ��[�U  1����  �tu /       Workout     �>\�U  @?\�U  �?\Some_stuffs_Some_stuffs_ �U  �B\�U  @C\�U   D\�U  �D\�U  ��Z��  O�u /      Meeting     `�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `[�U  z#[��  [�u /       Some_stuffs ��\�U  @�\�U  ��\justforfun_justforfun_ \�U  ��\�U  p�\�U  0�\�U  ��\�U  9]a��  �u /       Workout      �Y�U  �Y�U  0�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Y�U  -3���  �u /      Some_stuffs ��Y�U  ��Y�U  �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `�Y�U  (���  ��u /       Some_stuffs ��Y�U  ��Y�U  p�Yjustforfun_justforfun_ Y�U  ��Y�U  @�Y�U  ��Y�U  ��Y�U  �:���  :�u /      Birthday    p�Z�U  0�Z�U  ��Zjustforfun_justforfun_ Z�U  ��Z�U  ��Z�U  p�Z�U  ��Z�U  ��"��  v /       Appointment 0MZ�U  �MZ�U  pNZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   TZ�U  H����  �5v /       Appointment �%Y�U  �&Y�U  )YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �5Y�U  up���  �7v /      Appointment `�Z�U  �Z�U  `�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �Z�U  B\���  (8v /       Workout     ��Z�U  p�Z�U  0�ZSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ��Z�U  e�U��  �[v /      Birthday U  ��Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_ �U   �Z�U  ��Z�U   �Z�U  ��Z�U  h�c��  1_v /       Appointment �Z�U  �Z�U  `ZSome_stuffs_Some_stuffs_ �U  �Z�U  @Z�U    Z�U  � Z�U  D:���  �v /      Appointment 0�Z�U  ��Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�Z�U  tB���  �v /      Workout      [�U  �[�U  `[Some_stuffs_Some_stuffs_ �U   [�U  �[�U  `	[�U   
[�U  �.2��  ��v /       Workout     �r\�U  @s\�U   t\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   x\�U  ����  1�v /      Some_stuffs ��[�U  0�[�U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p�[�U  ��L��  �w /       Some_stuffs @�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_ �U  ��Z�U  `�Z�U   �Z�U  ��Z�U  pAN��  Fw /       Workout     0�[�U  ��[�U  p�[Some_stuffs_Some_stuffs_ �U  ��[�U  ��[�U  0�[�U  ��[�U  �E���  lDw /       Workout     ��Y�U  `�Y�U   �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  g���  
Hw /       Meeting     p;[�U  �;[�U  �<[This_stuffs_This_stuffs_ �U  p?[�U  �?[�U  p@[�U  �@[�U  D����  ,Kw /      Appointment �QZ�U  �RZ�U  �HZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �MZ�U  �	���  �nw /      Some_stuffs                    justforfun_justforfun_                                       ��#��  x�w /       Workout     ��[�U  P�[�U  �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��[�U  	(��  ��w /       Meeting     �Y[�U  pZ[�U  0[[This_stuffs_This_stuffs_ �U  �][�U  p^[�U  0_[�U  �_[�U  �c.��  0�w /      Appointment  _Z�U  �_Z�U  �`ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �eZ�U  f���  C�w /      Birthday                       justforfun_justforfun_                                       Y���  '�w /       Birthday    @�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_ �U  @�Z�U  ��Z�U  ��Z�U  @�Z�U  (pK��  )�w /       Meeting  nt p)]�U  �)]�U  p*]Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  @.]�U  �����  0x /       Meeting     ��Z�U  0�Z�U  ��Zjustforfun_justforfun_ _ his_stuffs_This_stuffs_ �U   �Z�U  �����  �x /       Appointment  �Y�U  ��Y�U  ��YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @�Y�U  ,�|��  M0x /      Workout �U  �<\�U  �=\�U  �_\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   B\�U  ZG���  �3x /       Birthday    �J\�U  PK\�U  L\justforfun_justforfun_ \�U  PN\�U  �N\�U  �O\�U  PP\�U  �2���  �5x /       Workout     �[�U  ��[�U  p�[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P�[�U  ؖ��   7x /       Appointment ��\�U  @�\�U  ��\Some_stuffs_Some_stuffs_ �U   �\�U  ��\�U   �\�U  ��\�U  �s)��  �\x /      Appointment @�[�U  ��[�U  @�[justforfun_justforfun_ _ �U  ��[�U  @�[�U   �[�U  ��[�U  X?1��  �^x /       Birthday                       This_stuffs_This_stuffs_                                     t{���  �|x /      Appointment ��X�U  @�X�U   YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �	Y�U  �����  �|x /       Meeting     PZ\�U  [\�U  �[\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��\�U  )���  ��x /       Some_stuffs �J^�U  PK^�U  �K^justforfun_justforfun_ ^�U  N^�U  �N^�U  O^�U  �O^�U  ��>��  ��x /       Workout     0TY�U   VY�U  @YYjustforfun_justforfun_ Y�U  paY�U  0bY�U  �eY�U  `fY�U  �@��  
�x /       Birthday     �]�U  ��]�U   �]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��]�U  
�F��  ��x /       Some_stuffs 0�\�U  ��\�U  0�\This_stuffs_This_stuffs_ �U  0]�U  �]�U  p]�U  0]�U  3�G��  ޥx /       Appointment p`[�U  �`[�U  �a[This_stuffs_This_stuffs_ �U  @d[�U  �d[�U  �e[�U   f[�U  �VT��  �x /       Some_stuffs  [�U  �[�U  `	[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �[�U  ����  �x /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �����  Y�x /       Some_stuffs ��Y�U  ��Y�U   �YThis_stuffs_This_stuffs_ �U  ��Y�U  ��Y�U   �Y�U  ��Y�U  �\|��  ��x /      Birthday fs ��\�U   �\�U  ��\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��\�U  <� ��  �y /      Some_stuffs EY�U  �EY�U  �HYjustforfun_justforfun_ Y�U  �PY�U  @QY�U  0TY�U   VY�U  I�(��  � y /       Appointment ��Z�U  ��Z�U  @�Zjustforfun_justforfun_ Z�U  @�Z�U   �Z�U  ��Z�U  ��Z�U  �̥��  �@y /       Birthday    ��Z�U  p�Z�U  0�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  ��;��  kgy /       Meeting �U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  B.[��  hoy /       Workout     �PY�U  @QY�U  0TYThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0bY�U  ��[��  �oy /      Meeting                        Some_stuffs_Some_stuffs_                                     �����  D�y /       Some_stuffs pO[�U  �O[�U  pP[This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  �T[�U  �����  N�y /       Appointment �v\�U   w\�U  �w\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �{\�U  ڀ���  w�y /       Appointment @k[�U  �k[�U  �l[This_stuffs_This_stuffs_ �U   o[�U  �o[�U  @p[�U   q[�U  �4���  (�y /      Workout                        justforfun_justforfun_                                       ّ���  �y /       Some_stuffs  Z�U  �Z�U  �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  pZ�U  i�r��  �y /       Birthday    �eY�U  `fY�U  �iYSome_stuffs_Some_stuffs_ �U  �sY�U  `tY�U  xY�U  �xY�U  �w��  �y /      Workout     ��\�U  ��\�U  0�\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�\�U  z���  ��y /       Birthday    �#[�U  p8[�U  p%[Some_stuffs_Some_stuffs_ �U  �'[�U  p([�U  0)[�U  �)[�U  �u���  Ļy /       Some_stuffs `�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  p�*�  e� /       Some_stuffs �Z�U  �Z�U  `ZThis_stuffs_This_stuffs_ �U  `Z�U  �Z�U  �Z�U  �%Z�U  ��A�  �j� /      Some_stuffs  �]�U  ��]�U  `�]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �]�U  �<��  ��� /       Birthday    �]�U  0]�U  �]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ]�U  e���  ��� /      Meeting     ��]�U  �]�U  ��]justforfun_justforfun_ ^�U  �^�U  ^�U  �^�U  ^�U  I_�  ��� /       Meeting ent @�[�U  ��[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �[�U  t�m�  ʷ� /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ����  �ۄ /      Appointment �e[�U   f[�U  �f[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �j[�U  ���  #�� /       Meeting     0�Z�U  �Z�U  p�Zjustforfun_justforfun_ Z�U  �Z�U  ��Z�U  0�Z�U  �Z�U  4���  b� /      Meeting �U  ��Z�U  `�Z�U   �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Z�U  4�%�  b(� /      Meeting     �[�U  P[�U  �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �[�U  ys-�  [*� /       Meeting     �y^�U  `z^�U  �z^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �~^�U  ����  �Q� /       Meeting     p^�U  �^�U  p^This_stuffs_This_stuffs_ �U  �^�U  � ^�U  p!^�U  0"^�U  ����  �S� /      Some_stuffs 0�Z�U  �Z�U  ��Zjustforfun_justforfun_ Z�U  @�Z�U  ��Z�U  �Z�U  p�Z�U  ��`	�  y� /       Appointment �Z�U  �Z�U  `Zjustforfun_justforfun_ Z�U  �Z�U  @Z�U    Z�U  � Z�U  ��e	�  Pz� /       Workout                        This_stuffs_This_stuffs_                                     @ g	�  �z� /       Some_stuffs                    Some_stuffs_Some_stuffs_                                     �Xl	�  �{� /      Workout �U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  ���	�  %�� /       Birthday    ��Z�U  `�Z�U   �Zjustforfun_justforfun_ Z�U  `�Z�U  ��Z�U  ��Z�U  `�Z�U  �-
�  ��� /      Some_stuffs ��Z�U  ��Z�U  `�Zjustforfun_justforfun_ Z�U   �Z�U  ��Z�U  `�Z�U   �Z�U  j�
�  Q�� /       Some_stuffs �H]�U  `I]�U  �I]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �M]�U  t��
�  �ƅ /      Birthday    �[�U  `[�U   [This_stuffs_This_stuffs_ �U  �[�U  `[�U   [�U  �[�U  ri�
�  Fǅ /       Birthday    �+Z�U  �,Z�U  �5ZThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  p1Z�U  ���
�  ZɅ /       Appointment ��Y�U  ��Y�U  P�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  Dt&�  ,� /      Workout     ��\�U   �\�U  ��\justforfun_justforfun_ \�U  P�\�U  Щ\�U  p�\�U  0�\�U  I,��  �� /       Workout     �[�U  ��[�U  p�[justforfun_justforfun_ [�U  ��[�U  �[�U  ��[�U  P�[�U  .ֽ�  �� /      Birthday    1]�U  �1]�U  @2]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �5]�U  ����  �� /       Meeting     ��Y�U  ��Y�U  `�Yjustforfun_justforfun_ Y�U  ��Y�U  ��Y�U  p�Y�U  0�Y�U  TK�  8� /       Some_stuffs 0:[�U  �:[�U  p;[Some_stuffs_Some_stuffs_ �U  �=[�U  �>[�U  p?[�U  �?[�U  K�K�  =8� /       Appointment P�[�U  �[�U  н[This_stuffs_This_stuffs_ �U  ��[�U  �[�U  ��[�U  P�[�U  9cQ�  �9� /       Birthday    �Z�U  ��Z�U   �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Z�U  ͰU�  �:� /       Meeting     P4\�U  �4\�U  P5\Some_stuffs_Some_stuffs_ �U  �7\�U  P8\�U  �8\�U  �9\�U  ��W�  N;� /       Meeting     �fZ�U  0rZ�U  �gZThis_stuffs_This_stuffs_ �U  �jZ�U  pkZ�U  0lZ�U  �lZ�U  ��[�  i<� /      Meeting ffs ��X�U  ��X�U  0�XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @�X�U  y{��  [_� /       Workout     @�\�U  ��\�U  @�\justforfun_justforfun_ \�U  ��\�U  ��\�U   �\�U  ��\�U  j���  �`� /       Some_stuffs ��\�U  ��\�U  @�\This_stuffs_This_stuffs_ �U  ��\�U   �\�U  ��\�U   �\�U  ���  ub� /       Meeting     ��X�U  @�X�U   YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �	Y�U  5��   c� /       Some_stuffs 0�\�U  ��\�U  ��\Some_stuffs_Some_stuffs_ �U  ��\�U  p�\�U  0�\�U  ��\�U  a�  Jh� /       Birthday    �&^�U  �'^�U   (^justforfun_justforfun_ _ �U   *^�U  �*^�U   +^�U  �+^�U  �͗�  C�� /       Meeting      �Z�U  ��Z�U  `�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   [�U  rP�  ��� /       Some_stuffs �]�U  @]�U  �]justforfun_justforfun_ ]�U  0!]�U  �!]�U  0"]�U  �"]�U  ��  ^�� /      Some_stuffs 5Y�U  �5Y�U  P8YSome_stuffs_Some_stuffs_ �U  @?Y�U  AY�U  EY�U  �EY�U  ��5�  ��� /       Meeting     ��Z�U  ��Z�U  p�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �Z�U  ���  :Ն /       Workout     �[�U  �[�U  [Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  [�U  LG��  �׆ /      Workout     `�Z�U   �Z�U  ��Zjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  `�Z�U  �:��  a؆ /       Workout     �Q[�U  pR[�U  0S[This_stuffs_This_stuffs_ �U  �U[�U  0V[�U  �V[�U  �W[�U  ���  �چ /       Appointment  �Z�U  ��Z�U   �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  �7��  �چ /       Workout     �Z�U  `�Z�U  �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P�Z�U  L�L�  !�� /      Meeting     ��X�U  ��X�U  0�XThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @�X�U  �L��  �"� /       Appointment �J\�U  PK\�U  L\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  PP\�U  ����  �'� /       Workout �U  ��]�U  ��]�U  �]justforfun_justforfun_ ]�U  ��]�U  P�]�U   �]�U  ��]�U  S��  �)� /      Workout     0iZ�U  �iZ�U  �jZSome_stuffs_Some_stuffs_ �U  pmZ�U  0nZ�U  �nZ�U  �oZ�U  z�~�  {K� /       Workout     �_\�U  `\�U  �>\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @C\�U  W��  `L� /       Appointment 0~[�U  �~[�U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0�[�U  �b��  cL� /       Birthday    �E[�U  0F[�U  �F[Some_stuffs_Some_stuffs_ �U  �I[�U  pJ[�U  0K[�U  �K[�U  䲒�  �P� /      Appointment xY�U  �xY�U  �|YSome_stuffs_Some_stuffs_ �U  ��Y�U  ��Y�U  p�Y�U  0�Y�U  U��  q� /      Workout     �a[�U  0b[�U  Pz[justforfun_justforfun_ [�U  �e[�U   f[�U  �f[�U  @g[�U  (��  �r� /       Meeting �U  �iY�U  �jY�U  @oYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P}Y�U  A���  ș� /       Some_stuffs p:^�U   ;^�U  �;^Some_stuffs_Some_stuffs_ �U  �=^�U  P>^�U  �>^�U  �?^�U  �:��  >�� /      Birthday     �Y�U  �Y�U  0�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Y�U  �G�  y�� /      Birthday    p3Z�U  04Z�U  �4Zjustforfun_justforfun_ Z�U  P8Z�U  9Z�U  �9Z�U  P:Z�U  Q.J�  �� /       Workout ent 0�]�U  �]�U  p�]Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  �]�U  !���  �� /       Meeting ffs @�]�U  ��]�U  ��]This_stuffs_This_stuffs_ �U  ��]�U  p�]�U  �]�U  Х]�U  ����  g� /      Meeting     @�Z�U  ��Z�U  �ZSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  p�Z�U  �1u�  �� /      Some_stuffs `�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_ �U  ��Z�U  `�Z�U   �Z�U  ��Z�U  [�{�  G� /       Birthday    ��[�U  ��[�U  @�[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��[�U  ��  j� /       Appointment xY�U  �xY�U  �|Yjustforfun_justforfun_ _ �U  ��Y�U  ��Y�U  p�Y�U  0�Y�U  �ؕ�  �� /       Appointment @j]�U   k]�U  �k]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �o]�U  -�  �8� /       Birthday    �<Z�U  P=Z�U  >ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  PCZ�U  d%�   9� /      Some_stuffs ��Z�U  ` [�U  `[This_stuffs_This_stuffs_ �U   [�U  �[�U  `[�U   [�U  ���  �[� /       Workout �U  ��]�U  `�]�U  ��]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �]�U  ����  �^� /      Meeting      �Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   �Z�U  �O�  �� /       Workout     �Y�U  `Y�U  �YSome_stuffs_Some_stuffs_ �U  �"Y�U  `#Y�U  �%Y�U  �&Y�U  �YT�  H�� /      Meeting     0_[�U  �_[�U  p`[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �d[�U  M��  �� /      Birthday    �.[�U  p/[�U  �/[justforfun_justforfun_ [�U  �2[�U  03[�U  �3[�U  p4[�U  ����  쫈 /       Meeting     �eY�U  `fY�U  �iYSome_stuffs_Some_stuffs_ �U  �sY�U  `tY�U  xY�U  �xY�U  �9��  k�� /       Meeting     �Z�U  �%Z�U  �Zjustforfun_justforfun_ Z�U  �!Z�U  @"Z�U   #Z�U  �#Z�U  �l��  x�� /       Meeting     )Z�U  �)Z�U  P*Zjustforfun_justforfun_ Z�U  �5Z�U  P6Z�U  �-Z�U  �.Z�U  �e��  ı� /       Appointment ��[�U  0�[�U  ��[Some_stuffs_Some_stuffs_ �U  0�[�U  �[�U  ��[�U  0�[�U  �m��  �؈ /      Meeting                        This_stuffs_This_stuffs_                                     �e�@�  �� /      Appointment 5Y�U  �5Y�U  P8Yjustforfun_justforfun_ Y�U  @?Y�U  AY�U  EY�U  �EY�U  zgA�  �Г /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             r�tA�  &ԓ /       Appointment `[�U   [�U  �[justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  `[�U  �-uA�  Eԓ /       Birthday    p�\�U  0�\�U  ��\Some_stuffs_Some_stuffs_ �U  p�\�U  ��\�U  p�\�U  ��\�U  i�yA�  qՓ /       Appointment ��X�U  @�X�U   Yjustforfun_justforfun_ Y�U  PY�U  Y�U   	Y�U  �	Y�U  ���A�  o�� /       Workout     @�\�U  P�\�U  ��\Some_stuffs_Some_stuffs_ �U  ��\�U  @�\�U  ��\�U  ��\�U  ���A�  E�� /       Appointment ��[�U  p�[�U  0�[Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ��[�U  EB�  ��� /      Meeting     �%]�U  p&]�U  �&]This_stuffs_This_stuffs_ �U  p)]�U  �)]�U  p*]�U   +]�U  (}B�  I�� /       Workout     �Z�U  ��Z�U   �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Z�U  |P�B�  � /      Appointment  �Z�U  ��Z�U  `�ZThis_stuffs_This_stuffs_ �U  ��Z�U  `�Z�U   �Z�U  �Z�U  �ʡB�  :!� /       Appointment p|Z�U  �|Z�U  �~ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  ���C�  �j� /      Meeting     @VZ�U   WZ�U  �WZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  pgZ�U  	��C�  �j� /       Some_stuffs ��Z�U  ��Z�U  0�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0�Z�U  �1TD�  o�� /      Some_stuffs pm^�U  �m^�U  pn^justforfun_justforfun_ ^�U  �p^�U  @q^�U  �q^�U  @r^�U  (WD�  )�� /       Birthday    @�[�U  ��[�U  ��[justforfun_justforfun_ [�U  @�[�U  ��[�U  @�[�U   �[�U   1�D�  ��� /       Meeting ent s[�U  �s[�U  t[This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  Px[�U  UQ�D�  ��� /      Appointment �\�U   \�U  �\This_stuffs_This_stuffs_ �U  `\�U   	\�U  �	\�U  �
\�U  ��E�  ��� /       Some_stuffs P[�U  [�U  �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �[�U  �x�E�  ��� /       Some_stuffs �v]�U  �w]�U   x]justforfun_justforfun_ ]�U  @z]�U  �z]�U  @{]�U   |]�U  ⇑E�  �� /       Appointment ��Z�U  `�Z�U   �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `�Z�U  �q�E�  �� /      Some_stuffs �Y�U  `Y�U  �Yjustforfun_justforfun_ _ �U  �Y�U   Y�U  �Y�U  @ Y�U  �%F�  �� /       Birthday    ��\�U  0�\�U  ��\Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  ��\�U  ��4F�  n� /       Workout     �+Z�U  �,Z�U  �5ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p1Z�U  *�7F�  I� /       Meeting     01[�U  �1[�U  �2[Some_stuffs_Some_stuffs_ �U  �4[�U  p5[�U  �5[�U  p6[�U  )P�F�  ).� /       Meeting     ��\�U  ��\�U  0�\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @�\�U  ���F�  75� /       Some_stuffs P'\�U  (\�U  �(\Some_stuffs_Some_stuffs_ �U  �+\�U  P,\�U  �,\�U  P-\�U  x�YG�  {V� /       Some_stuffs �[�U  0�[�U  ��[Some_stuffs_Some_stuffs_ �U  p�[�U  0�[�U  ��[�U  0�[�U  ��H�  E�� /      Meeting      B^�U  �B^�U   C^Some_stuffs_Some_stuffs_ �U  `E^�U  F^�U  �F^�U  G^�U  �H�  ��� /       Some_stuffs ��\�U  ��\�U  0�\Some_stuffs_Some_stuffs_ �U  ��\�U  @�\�U  ��\�U  @�\�U  ��H�  ã� /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             l�5I�  UЕ /      Appointment К]�U  P�]�U  Л]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��]�U  ��:I�  �ѕ /       Birthday    ��]�U  p�]�U  �]justforfun_justforfun_ _ �U  Ч]�U  P�]�U  Ш]�U  ��]�U  ��I�  �� /      Some_stuffs �[�U  ��[�U  p�[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P�[�U  ��I�  �� /       Meeting ffs �5Z�U  P6Z�U  �-ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �2Z�U  ���I�  �� /       Meeting     �[�U  ��[�U  ��[This_stuffs_This_stuffs_ �U  ��[�U  P�[�U  �[�U  ��[�U  ��I�  �� /       Appointment p^�U  �^�U  p^Some_stuffs_Some_stuffs_ �U  �^�U  � ^�U  p!^�U  0"^�U  �PYJ�  �� /       Meeting     �Z�U  �Z�U  `ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  � Z�U  M�jJ�  a� /      Meeting     �QZ�U  �RZ�U  �HZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �MZ�U  	�-L�  Ւ� /       Some_stuffs �[�U  0�[�U  ��[Some_stuffs_Some_stuffs_ �U  p�[�U  0�[�U  ��[�U  0�[�U  �U/L�  I�� /      Appointment  �Y�U  ЕY�U   �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  (I�L�  ɳ� /       Birthday    �$\�U  P%\�U  &\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  +\�U  �ڳL�  6�� /       Appointment 0[[�U  �[[�U  0\[This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  �`[�U  �~OM�  ݖ /       Birthday U  0�]�U  ��]�U  p�]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p�]�U  a,QM�  |ݖ /       Meeting      eZ�U  �eZ�U  �fZThis_stuffs_This_stuffs_ �U  0iZ�U  �iZ�U  �jZ�U  pkZ�U  �=TM�  Eޖ /      Workout  nt P^�U  �^�U  P^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0^�U  l
�M�  � /      Appointment  �Y�U  �Y�U  0�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Y�U  ��M�  � /       Birthday      Z�U  � Z�U  �!ZSome_stuffs_Some_stuffs_ �U  �$Z�U  p-Z�U  &Z�U  �&Z�U  ���N�  �+� /      Some_stuffs 0K[�U  �K[�U  c[justforfun_justforfun_ [�U  pO[�U  �O[�U  pP[�U  0Q[�U  ��O�  XR� /       Appointment  �Y�U  �Y�U  0�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Y�U  �&O�  �U� /       Appointment �
]�U  0]�U  �]Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  �]�U  ��-O�  rW� /      Workout     �Z�U  �Z�U  �ZSome_stuffs_Some_stuffs_ �U  0	Z�U  �	Z�U  p
Z�U  0Z�U  ���O�  �~� /       Meeting     `Z�U   Z�U  �Zjustforfun_justforfun_ Z�U  �Z�U  �%Z�U  �Z�U  @Z�U  ą�O�  � /      Birthday    �Z�U  �Z�U  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Z�U  ��HP�  ��� /       Appointment �(\�U  �)\�U  P*\This_stuffs_This_stuffs_ �U  �,\�U  P-\�U  .\�U  �.\�U  ��PP�  �� /       Appointment                    Some_stuffs_Some_stuffs_                                     �SP�  ʢ� /       Meeting     �\�U  p\�U  0\This_stuffs_This_stuffs_ �U  p\�U  �\�U  �\�U  p\�U  �@UP�  #�� /       Some_stuffs �PY�U  @QY�U  0TYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0bY�U  I��P�  �ŗ /       Birthday    ��X�U  @�X�U   YSome_stuffs_Some_stuffs_ �U  PY�U  Y�U   	Y�U  �	Y�U  4�P�  �ŗ /      Birthday U  ��Y�U  ��Y�U  p�YThis_stuffs_This_stuffs_ �U  ��Y�U  @�Y�U  ��Y�U  ��Y�U  :��P�  Ǘ /       Appointment  �Z�U  ��Z�U  `�ZThis_stuffs_This_stuffs_ �U  ��Z�U  ��Z�U  `�Z�U   �Z�U  ,K�P�  	ɗ /       Birthday    @�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_ �U  ��Z�U   �Z�U  ��Z�U  ��Z�U  sz�P�  �˗ /       Appointment �/[�U  p0[�U  01[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p5[�U  l�R�  5� /      Workout     p�Z�U  0�Z�U  ��ZSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  0�Z�U  )fR�  �� /       Some_stuffs 0]�U  �]�U  p]This_stuffs_This_stuffs_ �U  �]�U  0]�U  �]�U  0]�U  2R�R�  ><� /       Meeting     ��Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Z�U  DA�R�  L?� /      Birthday nt ��Z�U  ��Z�U  @�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  y��R�  ;B� /       Workout �U  ��Z�U  `�Z�U   �Zjustforfun_justforfun_ Z�U  ��Z�U  ��Z�U  0�Z�U  ��Z�U  ,l|�  �� /      Workout     ;Z�U  �;Z�U  �<ZThis_stuffs_This_stuffs_ �U  �?Z�U  �@Z�U  PAZ�U  �AZ�U  a�r|�  <� /       Some_stuffs ��\�U  p�\�U  0�\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p�\�U  �}�  �� /       Some_stuffs �<Z�U  P=Z�U  >ZSome_stuffs_Some_stuffs_ �U  PAZ�U  �AZ�U  �BZ�U  PCZ�U  ��}�  	8� /      Meeting     ppZ�U  0qZ�U  p}ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0vZ�U  �֘}�  �9� /       Meeting ffs `[�U   [�U  �[Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U   [�U  �H�}�  �;� /       Workout     �^�U  �^�U  `^This_stuffs_This_stuffs_ �U  �^�U  `^�U  �^�U  �^�U  0��}�  �>� /       Meeting �U  �Z�U  @Z�U  PZjustforfun_justforfun_ Z�U  PZ�U  �Z�U  �Z�U  PZ�U  �,~�  j_� /       Workout     �5[�U  p6[�U  07[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �:[�U  �C6~�  �a� /      Some_stuffs ��Y�U  `�Y�U   �YSome_stuffs_Some_stuffs_ �U  p�Y�U  0�Y�U  ��Y�U  ��Y�U  R�C~�  Re� /       Birthday    p"\�U  �"\�U  �#\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  (\�U   k�~�  4�� /       Some_stuffs ��Y�U  ��Y�U  p�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  ��~�  `�� /       Some_stuffs  �\�U  ��\�U  ��\justforfun_justforfun_ \�U  ��\�U  0�\�U  ��\�U  0�\�U  ���~�  b�� /       Appointment 0b]�U  �b]�U  pc]Some_stuffs_Some_stuffs_ �U  �e]�U  pf]�U  �f]�U  pg]�U  e�~�  ��� /       Appointment `�Z�U   �Z�U  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �Z�U  ���~�  :�� /      Meeting     p�Y�U  0�Y�U  0�Yjustforfun_justforfun_ Y�U   �Y�U  ��Y�U  ��Y�U  p�Y�U  �8o�  ��� /       Appointment  �[�U  ��[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��[�U  ��v�  볣 /       Meeting      �\�U  ��\�U   �\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �\�U  ����  �ң /       Appointment ��Z�U  0�Z�U  �ZSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ��Z�U  vM��  �ӣ /      Birthday    ��Z�U   �Z�U   �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `�Z�U  ���  �֣ /       Birthday    )Z�U  �)Z�U  P*ZThis_stuffs_This_stuffs_ �U  �5Z�U  P6Z�U  �-Z�U  �.Z�U  a���  \ۣ /       Birthday    P4\�U  �4\�U  P5\This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  �9\�U   C���  4�� /       Some_stuffs �;Y�U  `<Y�U  @?YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `MY�U  Kݎ��  ��� /       Meeting ffs ��\�U   �\�U  ��\This_stuffs_This_stuffs_ �U  ��\�U  @�\�U  ��\�U  @�\�U  �ꑀ�  e�� /       Meeting     ��\�U  0�\�U  �\Some_stuffs_Some_stuffs_ �U  p�\�U  �\�U  p�\�U  �\�U  hw���  ` � /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             i����  �� /       Workout      �Z�U  ��Z�U  `�ZThis_stuffs_This_stuffs_ �U  ��Z�U  ��Z�U  `�Z�U   �Z�U  I�0��  %� /       Meeting     �eY�U  `fY�U  �iYjustforfun_justforfun_ Y�U  �sY�U  `tY�U  xY�U  �xY�U  �}7��  �&� /      Appointment p�Y�U  0�Y�U  ��YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  �>��  �(� /       Some_stuffs                    justforfun_justforfun_                                       1�Ɂ�  >L� /       Some_stuffs 0�X�U  ��X�U  ��Xjustforfun_justforfun_ X�U  ��X�U  ��X�U  ��X�U  ��X�U  Dn΁�  lM� /      Meeting     `\�U  �\�U  `\This_stuffs_This_stuffs_ �U  �\�U   \�U  �\�U  `\�U  :�ρ�  �M� /       Some_stuffs ��]�U  @�]�U  ��]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��]�U  ��R��  Qo� /      Workout     �%Y�U  �&Y�U  )YSome_stuffs_Some_stuffs_ �U  �1Y�U  �2Y�U  5Y�U  �5Y�U  	%]��  �q� /       Birthday    �[�U  �[�U  `[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �$[�U  p��  ��� /       Some_stuffs ��Y�U  ��Y�U  p�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  }����  ߽� /      Birthday    ��X�U  ��X�U  0�XThis_stuffs_This_stuffs_ �U   �X�U  ��X�U  ��X�U  @�X�U  �酃�   /       Workout      �Y�U  ��Y�U  ��YThis_stuffs_This_stuffs_ �U  P�Y�U  �Y�U  ��Y�U  ��Y�U  2u���  �� /       Some_stuffs 0\�U  �\�U  0\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @>\�U  3!���  �ä /       Some_stuffs                    justforfun_justforfun_ _Some_stuffs_Some_stuffs_             �"��  � /       Workout     �8\�U  �9\�U  P:\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `\�U  ��4��  �� /      Appointment Pu[�U  �u[�U  Pv[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p�[�U  Ђ5��  �� /       Appointment ��X�U  ��X�U  0�XSome_stuffs_Some_stuffs_ �U   �X�U  ��X�U  ��X�U  @�X�U   nɄ�  �� /       Birthday    ��X�U  ��X�U  0�XThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @�X�U  ��ʄ�  $� /       Some_stuffs @�\�U  P�\�U  ��\This_stuffs_This_stuffs_ �U  ��\�U  @�\�U  ��\�U  ��\�U  kτ�  1� /       Some_stuffs �\�U  @>\�U  \justforfun_justforfun_ \�U  @!\�U  �!\�U  p"\�U  �"\�U  mф�  �� /      Workout �U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  40҄�  �� /       Workout     `�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `�Z�U  �Dc��  "8� /       Birthday    ��Y�U  ��Y�U  p�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  
�c��  58� /       Workout     ��X�U  ��X�U  0�XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @�X�U  �l��  �:� /      Birthday    �Z�U  p�Z�U  ��ZSome_stuffs_Some_stuffs_ �U  ��Z�U  p�Z�U  0�Z�U  ��Z�U  ����  �\� /      Birthday U  t[�U  �t[�U  Pu[Some_stuffs_Some_stuffs_ �U  �w[�U  Px[�U  �x[�U  �y[�U  kq���  q�� /       Some_stuffs �cZ�U  `dZ�U   eZSome_stuffs_Some_stuffs_ �U  �gZ�U  phZ�U  0iZ�U  �iZ�U  ^Ō��  K�� /      Meeting     �Y�U  `Y�U  �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `#Y�U  p���  f�� /       Appointment 0TY�U   VY�U  @YYThis_stuffs_This_stuffs_ �U  paY�U  0bY�U  �eY�U  `fY�U  �蕆�  ��� /       Some_stuffs �+Z�U  �,Z�U  �5ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p1Z�U  �l&��  ��� /       Workout     0�\�U  ��\�U  ��\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��\�U  ����  �Υ /      Some_stuffs  
^�U  �
^�U   ^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �^�U  x0���  {ҥ /       Meeting     �~Z�U  0Z�U  �ZThis_stuffs_This_stuffs_ �U  ��Z�U  ��Z�U  p�Z�U  0�Z�U  b!S��  ��� /       Some_stuffs ��[�U  P�[�U  ��[Some_stuffs_Some_stuffs_ �U  P�[�U  ��[�U  ��[�U  `�[�U  ��T��  �� /       Birthday nt  �]�U  ��]�U  0�]This_stuffs_This_stuffs_ �U   �]�U  ��]�U   �]�U  ��]�U  t�Z��  ��� /      Birthday                       Some_stuffs_Some_stuffs_                                     X���  �!� /       Some_stuffs P�Y�U  �Y�U  ��YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  �v���  �$� /       Workout      Z�U  �Z�U  �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  pZ�U  �2w��  aC� /       Meeting     p�Z�U  0�Z�U  ��Zjustforfun_justforfun_ _ �U  p�Z�U  0�Z�U   �Z�U  ��Z�U  Rِ��  �I� /       Meeting     �-]�U  @.]�U  �.]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �2]�U  5���  �J� /      Meeting     ppZ�U  0qZ�U  p}ZSome_stuffs_Some_stuffs_ �U  0tZ�U  �tZ�U  puZ�U  0vZ�U  ���  �m� /      Meeting     �EZ�U  PFZ�U  GZSome_stuffs_Some_stuffs_ �U  �HZ�U  �IZ�U  0JZ�U  �JZ�U  MN���  A�� /      Birthday U  P�^�U  �^�U  ��^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �^�U  �վ��  A�� /       Meeting ent p�[�U  0�[�U  ��[Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  �[�U  t����  j� /      Meeting     �9Z�U  P:Z�U  ;ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �@Z�U  ��z��  �� /      Meeting     @�Z�U  ��Z�U  �ZSome_stuffs_Some_stuffs_ �U  p�Z�U  ��Z�U  ��Z�U  p�Z�U  �p���  �� /       Some_stuffs �\�U  ��\�U  @�\justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  @�\�U  yr��  �/� /       Birthday fs P~^�U  �~^�U  P^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @�^�U  �j!��  �3� /      Workout     ��Z�U  0�Z�U  ��ZThis_stuffs_This_stuffs_ �U  `�Z�U  ��Z�U  `�Z�U   �Z�U  |DÍ�  �\� /      Workout ffs @�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �Z�U  �����  �*� /       Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �O���  X+� /       Some_stuffs �g\�U  0h\�U  �h\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �l\�U  ����  W� /       Workout �U  �HY�U  �IY�U  �LYjustforfun_justforfun_ Y�U  0TY�U   VY�U  @YY�U   ZY�U  �����  �X� /      Birthday    p�Y�U  0�Y�U  0�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�Y�U  ��-��  Nz� /       Meeting     `�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_ �U  `�Z�U   �Z�U  �Z�U  `�Z�U  ��7��  �|� /      Some_stuffs ��Y�U  p�Y�U  ��Yjustforfun_justforfun_ Y�U   �Y�U  �Y�U  0�Y�U  �Y�U  �'>��  �~� /       Some_stuffs 0b]�U  �b]�U  pc]Some_stuffs_Some_stuffs_ �U  �e]�U  pf]�U  �f]�U  pg]�U  �HA��  N� /       Some_stuffs ��[�U   �[�U  ��[Some_stuffs_Some_stuffs_ �U  ��[�U   �[�U  ��[�U  @�[�U  ��չ�  P�� /      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �F۹�  ��� /       Some_stuffs p�Z�U  ��Z�U  p�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�Z�U  <#\��  �ǲ /      Some_stuffs EY�U  �EY�U  �HYjustforfun_justforfun_ Y�U  �PY�U  @QY�U  0TY�U   VY�U  	���  �� /       Birthday U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  �0���  �� /       Some_stuffs  �X�U  ��X�U  ��XSome_stuffs_Some_stuffs_ �U  �Y�U  pY�U  PY�U  Y�U  �����  � /      Meeting     ��Y�U  ��Y�U  p�YThis_stuffs_This_stuffs_ �U  ��Y�U  @�Y�U   �Y�U  ��Y�U  {
��  ;�� /       Birthday nt �Z�U  `Z�U   ZSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  �Z�U  Û��  �� /       Meeting  fs �Z�U  ��Z�U  p�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �Z�U  |Ǩ��  �� /      Appointment                    This_stuffs_This_stuffs_                                     C0���  �d� /       Workout     ��^�U  �^�U  ��^justforfun_justforfun_ ^�U  ��^�U  @�^�U  ��^�U  @�^�U  �rμ�  h� /       Birthday    �PY�U  @QY�U  0TYSome_stuffs_Some_stuffs_ �U  P]Y�U  ^Y�U  paY�U  0bY�U  UҼ�  �h� /      Some_stuffs 0�Z�U  ��Z�U  ��Zjustforfun_justforfun_ Z�U  p�Z�U  ��Z�U  ��Z�U  0�Z�U  ��ܼ�  �k� /       Some_stuffs 0�\�U  ��\�U  p�\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P�\�U  �8c��  #�� /       Workout     0MZ�U  �MZ�U  pNZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   TZ�U  �1j��  쏳 /       Birthday    �p^�U  @q^�U  �q^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �u^�U  ��k��  Y�� /       Some_stuffs                    This_stuffs_This_stuffs_                                     Hg���  ݵ� /       Appointment P�Y�U  �Y�U  ��YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  ����  ��� /      Meeting     ��\�U   �\�U  ��\justforfun_justforfun_ \�U  p�\�U  ��\�U  ��\�U  @�\�U  T����  2س /       Appointment 0�\�U  ��\�U  0�\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0]�U  DN���  lٳ /      Some_stuffs ��Y�U  p�Y�U  ��YThis_stuffs_This_stuffs_ �U  �Y�U  ��Y�U   �Y�U  �Y�U  ����  �۳ /       Birthday    EY�U  �EY�U  �HYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   VY�U  �����  �ܳ /       Workout ffs �[�U  �[�U  `[This_stuffs_This_stuffs_ �U   [�U  �[�U  �[�U  �$[�U  N����  �ݳ /       Appointment �\�U  ��\�U   �\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �\�U  ���  ޳ /       Birthday U   �]�U  ��]�U   �]This_stuffs_This_stuffs_ �U   �]�U  ��]�U  `�]�U  ��]�U  �J���  �߳ /       Birthday    &\�U  �&\�U  P'\justforfun_justforfun_ \�U  P*\�U  +\�U  �+\�U  P,\�U  P+��  �� /       Meeting     �Y�U   Y�U  �YSome_stuffs_Some_stuffs_ �U  �%Y�U  �&Y�U  )Y�U  �)Y�U  �J+��  �� /       Birthday U  P�[�U  �[�U  й[This_stuffs_This_stuffs_ �U  P�[�U  �[�U  н[�U  ��[�U  b0��  � /       Some_stuffs P�[�U  ��[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `�[�U  �yƿ�  �*� /      Appointment @�[�U  ��[�U  @�[Some_stuffs_Some_stuffs_ �U  ��[�U  ��[�U   �[�U  ��[�U  #�ƿ�  �*� /       Meeting     �Q\�U  PR\�U  S\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  W\�U  ӿ�  �-� /       Appointment `�Y�U   �Y�U   �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  ��տ�  �.� /       Birthday    `�Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  =Q��  $N� /      Appointment                    justforfun_justforfun_                                       �D\��  �P� /       Birthday    0�Z�U  �Z�U  p�ZThis_stuffs_This_stuffs_ �U  �Z�U  ��Z�U  0�Z�U  �Z�U  �]��  VQ� /       Meeting     pf\�U  �f\�U  �g\justforfun_justforfun_ \�U   j\�U  �j\�U  @k\�U  �k\�U  ����  �t� /       Workout     `�Z�U   �Z�U  ��Zjustforfun_justforfun_ Z�U  `�Z�U   �Z�U  �Z�U  `�Z�U  &����  �w� /      Some_stuffs Pz[�U  �z[�U  @d[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �h[�U  `����  �z� /       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_              ����  ��� /       Meeting �U  ��Z�U  0�Z�U  �ZSome_stuffs_Some_stuffs_ �U  �Z�U  p�Z�U  ��Z�U  ��Z�U  �:���  ��� /       Some_stuffs ��\�U   �\�U  ��\justforfun_justforfun_ \�U  �\�U  ��\�U  �\�U  ��\�U  �{���  ��� /      Meeting �U  �[�U  �[�U  P[Some_stuffs_Some_stuffs_ �U  �[�U  �[�U   [�U  � [�U  ��"��  CŴ /       Some_stuffs                    Some_stuffs_Some_stuffs_                                     ��*��  aǴ /       Birthday    �?\�U  �@\�U  @A\Some_stuffs_Some_stuffs_ �U   D\�U  �D\�U  0E\�U  �E\�U  p],��  �Ǵ /       Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             v:��  J˴ /      Some_stuffs �+Z�U  �,Z�U  �5ZThis_stuffs_This_stuffs_ �U  0/Z�U  �/Z�U  �0Z�U  p1Z�U  `����  �� /       Some_stuffs �F[�U  �G[�U  pH[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �c[�U  a����  �� /       Some_stuffs  	Y�U  �	Y�U  �YSome_stuffs_Some_stuffs_ �U  �Y�U  `Y�U  �Y�U  `Y�U  �����  g� /      Some_stuffs �K^�U  PL^�U  �L^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �P^�U  �_���  �� /       Meeting      �Z�U  ��Z�U  0�ZSome_stuffs_Some_stuffs_ �U  0�Z�U  ��Z�U  p�Z�U  ��Z�U  mT��  u� /      Appointment p�Z�U  0�Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0�Z�U  ��^��  8� /       Meeting     �[�U  [�U  �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  #[�U  ����  �7� /      Meeting     P4\�U  �4\�U  P5\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �9\�U  �C���  0e� /       Meeting     �Z�U  pZ�U  0	Zjustforfun_justforfun_ Z�U  �Z�U  �Z�U  �Z�U  @Z�U  d:��  @�� /      Appointment p�Z�U  0�Z�U  ��ZThis_stuffs_This_stuffs_ �U  0�Z�U  �Z�U  ��Z�U  0�Z�U  �((��  N�� /       Workout     ��Y�U  ��Y�U  P�YThis_stuffs_This_stuffs_ �U  �Y�U  ��Y�U  0�Y�U  ��Y�U  �,5��  ��� /       Appointment �H\�U  PI\�U  �I\justforfun_justforfun_ _ �U  L\�U  �L\�U  PM\�U  �M\�U  I����  }�� /       Birthday                       This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_             �����  1�� /      Some_stuffs 0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  "����  ��� /       Some_stuffs �%Y�U  �&Y�U  )YSome_stuffs_Some_stuffs_ �U  �1Y�U  �2Y�U  5Y�U  �5Y�U  �#F��  �Ե /       Birthday    EY�U  �EY�U  �HYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   VY�U  �!a��  m۵ /       Birthday nt �l]�U  @m]�U  �m]Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  �q]�U  m�b��  �۵ /      Meeting �U  �#[�U  p8[�U  p%[Some_stuffs_Some_stuffs_ �U  �'[�U  p([�U  0)[�U  �)[�U  �����  F� /      Birthday nt ��]�U  @�]�U  ��]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P�]�U  @Zx��  �"� /       Birthday U  ��\�U  @�\�U  ��\This_stuffs_This_stuffs_ �U  ��\�U  @�\�U  ��\�U  ��\�U  �az��  m#� /       Meeting     �V^�U   W^�U  �W^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p[^�U  �;���  �%� /      Appointment P�^�U  ��^�U  P�^Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   �^�U  Ѿ���  b(� /       Appointment @ \�U  � \�U  @!\This_stuffs_This_stuffs_ �U  �#\�U  P$\�U  �$\�U  P%\�U  ����  �*� /       Meeting ffs ��Y�U  ��Y�U  p�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  �G��  \L� /      Workout     �8[�U  p9[�U  0:[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �>[�U   ?���  �p� /       Some_stuffs P�Y�U  �Y�U  ��YThis_stuffs_This_stuffs_ �U   �Y�U  ��Y�U  ��Y�U  ��Y�U  �ͩ��  q� /      Appointment @}\�U  �}\�U  @~\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �\�U  �Ѵ��  �s� /       Appointment �Z�U  p�Z�U  ��Zjustforfun_justforfun_ Z�U  ��Z�U  p�Z�U  0�Z�U  ��Z�U  ��A��  �� /       Birthday fs �F[�U  �G[�U  pH[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �c[�U  HG��  ]�� /       Meeting ent ��Y�U  ��Y�U  �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `�Y�U  >V��  ?�� /       Appointment                    This_stuffs_This_stuffs_                                     T�W��  ��� /       Meeting     ��\�U  @�\�U  ��\This_stuffs_This_stuffs_ �U   �\�U  ��\�U  @�\�U  ��\�U  ]+a��  �� /      Birthday     [�U  �[�U  `	[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �[�U  ^���  ��� /       Some_stuffs                    Some_stuffs_Some_stuffs_                                     �����  �¶ /       Birthday    P[�U  [�U  �[This_stuffs_This_stuffs_ �U   [�U  � [�U  P![�U  "[�U  1����  ^ƶ /       Birthday nt ��Y�U  `�Y�U   �YSome_stuffs_Some_stuffs_ �U  p�Y�U  0�Y�U  ��Y�U  ��Y�U  ͌�p,�  Q2 &/      Some_stuffs p\�U  �\�U  �\justforfun_justforfun_ \�U  \�U  �\�U  @ \�U  � \�U  Zp�p,�  '7 &/       Birthday    �D]�U  E]�U  �E]justforfun_justforfun_ ]�U  �G]�U  0H]�U  �H]�U  `I]�U  (��p,�  �7 &/       Meeting     �Z�U  pZ�U  0	ZSome_stuffs_Some_stuffs_ �U  �Z�U  �Z�U  �Z�U  @Z�U  ��iq,�  �\ &/      Workout     @SZ�U   TZ�U  �TZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �YZ�U  ��tq,�  d_ &/       Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             -vq,�  �_ &/       Some_stuffs �/[�U  p0[�U  01[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p5[�U  �׀q,�  �b &/       Some_stuffs ��Z�U  ��Z�U  @�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Z�U  ���q,�  �� &/       Birthday nt @�[�U  ��[�U  ��[justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  P�[�U  ��r,�  � &/       Birthday nt ��Z�U  p�Z�U  0�Zjustforfun_justforfun_ _This_stuffs_This_stuffs_ �U  ��Z�U  Yץr,�  �� &/       Some_stuffs �Z�U  ��Z�U  @�ZSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  ��Z�U  ��r,�  � &/      Birthday    �Z�U  �Z�U  `ZThis_stuffs_This_stuffs_ �U  �Z�U  @Z�U    Z�U  � Z�U  �Ьr,�  P� &/       Birthday    �;\�U  P<\�U  �<\This_stuffs_This_stuffs_ �U  �>\�U  @?\�U  �?\�U  �@\�U  �z+s,�  �� &/      Some_stuffs @v^�U  �v^�U  �w^This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  `{^�U  �Ds,�  � &/       Meeting     P[�U  [�U  �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �[�U  ���s,�  I� &/      Workout �U  ��^�U   �^�U  ��^This_stuffs_This_stuffs_ �U  ��^�U  0�^�U  ��^�U  0�^�U  q�s,�  &� &/       Workout     &\�U  �&\�U  P'\This_stuffs_This_stuffs_ �U  P*\�U  +\�U  �+\�U  P,\�U  Tsut,�  6$&/      Meeting ent   Z�U  � Z�U  �!ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �&Z�U  D!u,�  LK&/      Birthday     �Z�U  ��Z�U  0�ZThis_stuffs_This_stuffs_ �U  0�Z�U  ��Z�U  p�Z�U  ��Z�U  �	�u,�  �k&/      Workout     @�\�U  ��\�U  p�\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  Н\�U  *z�u,�  il&/       Birthday    pH[�U  0I[�U  �I[This_stuffs_This_stuffs_ �U  c[�U  �c[�U  N[�U  �N[�U  �M�u,�  �n&/       Some_stuffs                    justforfun_justforfun_                                       9��u,�  Sr&/       Workout �U  p�\�U  �\�U  p�\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��\�U  �=6v,�  �&/       Meeting     puZ�U  0vZ�U  �vZSome_stuffs_Some_stuffs_ �U  �yZ�U  0zZ�U  �zZ�U  �{Z�U   <v,�  ��&/       Birthday    �%Y�U  �&Y�U  )YSome_stuffs_Some_stuffs_ �U  �1Y�U  �2Y�U  5Y�U  �5Y�U  2�=v,�  ��&/       Workout ffs  eZ�U  �eZ�U  �fZThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  pkZ�U  ��v,�  +�&/       Birthday    �/[�U  p0[�U  01[justforfun_justforfun_ _ �U  �3[�U  p4[�U  �4[�U  p5[�U  <l�v,�  W�&/      Workout �U  0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  ���v,�  x�&/       Appointment 0�\�U  ��\�U  ��\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��\�U  �Mdw,�  n�&/       Meeting                        This_stuffs_This_stuffs_                                     �N�w,�  �	&/       Some_stuffs Ш]�U  ��]�U   �]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��]�U  |��w,�  _
&/      Meeting �U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��X�U  q��w,�  f&/       Appointment p�Z�U  0�Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0�Z�U  䲍x,�  �0&/      Workout                        This_stuffs_This_stuffs_                                     ��!y,�  �V&/       Appointment �o\�U  �p\�U  @q\This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U   v\�U  �y8y,�  H\&/      Meeting                        This_stuffs_This_stuffs_                                     X½y,�  g~&/       Birthday                       justforfun_justforfun_                                       2i�y,�  ��&/       Appointment �\Z�U   ]Z�U  @SZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @XZ�U  UU�y,�  v�&/      Appointment `	[�U   
[�U  �
[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `[�U  1�Xz,�  �&/       Meeting     �p^�U  @q^�U  �q^justforfun_justforfun_ ^�U  �s^�U  �t^�U  @u^�U  �u^�U  ��]z,�  c�&/       Some_stuffs �k]�U  @l]�U  �l]This_stuffs_This_stuffs_ �U   o]�U  �o]�U  @p]�U  �p]�U  ���z,�  3�&/      Birthday    @�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @�Z�U  H��{,�  }�&/       Meeting     `Z�U   Z�U  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @Z�U  *B|,�  i&/       Some_stuffs �l[�U   m[�U  �m[This_stuffs_This_stuffs_ �U  @p[�U   q[�U  �q[�U  Pr[�U  )�|,�  �&/       Appointment PAZ�U  �AZ�U  �BZThis_stuffs_This_stuffs_ �U  �EZ�U  PFZ�U  GZ�U  �GZ�U  <�0|,�  �&/      Meeting �U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  *#�|,�  	@&/       Workout     @oY�U   pY�U  �sYjustforfun_justforfun_ Y�U  �|Y�U  P}Y�U   �Y�U  ��Y�U  d=�|,�  B&/       Meeting     �%Y�U  �&Y�U  )YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �5Y�U  ��|,�  �F&/      Meeting     7Z�U  �7Z�U  P8ZSome_stuffs_Some_stuffs_ �U  ;Z�U  �;Z�U  �<Z�U  P=Z�U  S�|,�  2G&/       Workout     �fZ�U  0rZ�U  �gZThis_stuffs_This_stuffs_ �U  �jZ�U  pkZ�U  0lZ�U  �lZ�U  �*�|,�  6G&/       Workout     07[�U  �7[�U  �L[This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  �;[�U  !�I},�  �f&/       Meeting                        Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_             �R},�  �h&/      Appointment p�Y�U  0�Y�U  0�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�Y�U  KQ^},�  l&/       Birthday nt �nZ�U  �oZ�U  ppZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �tZ�U  ��_},�  �l&/       Birthday nt  �^�U  ��^�U   �^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��^�U  `��~,�  |�&/       Appointment ��\�U   �\�U  ��\justforfun_justforfun_ \�U  p�\�U  0�\�U  ��\�U  0�\�U  l/,�  5�&/      Birthday fs 0�Z�U  ��Z�U  ��ZThis_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  p�Z�U  ���,�  �&/      Workout      �Y�U  ��Y�U  ��YThis_stuffs_This_stuffs_ �U  �Z�U  `Z�U   Z�U  �Z�U  ��,�  �&/       Some_stuffs  ;]�U  �;]�U  �<]This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  `@]�U  Ӊ�,�  B&/       Workout     �\�U  ��\�U   �\justforfun_justforfun_ _ �U   �\�U  ��\�U   �\�U  �\�U  �ּ,�  b&/       Meeting     `�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �Z�U  `0�,�  �&/       Birthday    P�Y�U  �Y�U  ��YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  ��Y�,�  �/&/      Appointment �Z�U  PZ�U  ZThis_stuffs_This_stuffs_ �U  `Z�U   Z�U  �Z�U  �Z�U  мg�,�  "3&/       Birthday     �Y�U  �Y�U  0�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Y�U  q��,�  fS&/       Workout     `�Z�U   �Z�U  ��Zjustforfun_justforfun_ Z�U  `�Z�U   �Z�U  ��Z�U  `�Z�U  �G��,�  ^W&/      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ��$�,�  �&/      Workout     �Y�U  `Y�U  �YSome_stuffs_Some_stuffs_ �U  �"Y�U  `#Y�U  �%Y�U  �&Y�U  ���,�  .�&/       Birthday    �Z�U  PZ�U  ZThis_stuffs_This_stuffs_ �U  `Z�U   Z�U  �Z�U  �Z�U  􉯂,�  ��&/       Workout     )Z�U  �)Z�U  P*ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �.Z�U  �ᰂ,�  ��&/       Birthday fs p�\�U  �\�U  p�\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��\�U  4��,�  �&/      Birthday U  xY�U  �xY�U  �|Yjustforfun_justforfun_ Y�U  ��Y�U  ��Y�U  p�Y�U  0�Y�U  ꨱ�,�  !�&/       Some_stuffs pNZ�U  0OZ�U  �OZThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  �UZ�U  %���,�  ��&/       Some_stuffs @i[�U  �i[�U  @j[justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  �n[�U  ��g�,�  �v&/      Appointment ��Z�U  p�Z�U  0�Zjustforfun_justforfun_ Z�U  ��Z�U  p�Z�U  0�Z�U  ��Z�U  ��~�,�  �|&/       Workout �U  pf\�U  �f\�U  �g\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �k\�U  �g�,�  V�&/       Meeting     �+Z�U  �,Z�U  �5Zjustforfun_justforfun_ Z�U  0/Z�U  �/Z�U  �0Z�U  p1Z�U  e�,�  ��&/      Birthday    �6]�U   7]�U  �7]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �;]�U  YP�,�  '�&/       Appointment ��Z�U  p�Z�U  0�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �Z�U  K��,�  ��&/      Appointment �F[�U  �G[�U  pH[justforfun_justforfun_ [�U  0K[�U  �K[�U  c[�U  �c[�U  ���,�  ,�&/       Some_stuffs �Z�U  �%Z�U  �Zjustforfun_justforfun_ _ �U  �!Z�U  @"Z�U   #Z�U  �#Z�U  �秭,�  ��&/       Some_stuffs �m[�U  �n[�U   o[justforfun_justforfun_ _ �U  �q[�U  Pr[�U  s[�U  �s[�U  Ji��,�  �&/       Workout     ��\�U   �\�U  ��\This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  `�\�U  |/9�,�  ��&/      Meeting ffs �Z�U  p�Z�U  ��ZThis_stuffs_This_stuffs_ �U  ��Z�U  p�Z�U  0�Z�U  ��Z�U  ,AѮ,�  �&/      Birthday     �Y�U  �Y�U  0�Yjustforfun_justforfun_ Y�U  ��Y�U  ��Y�U  P�Y�U  �Y�U  	`Ѯ,�  �&/       Appointment `]�U   ]�U  �]justforfun_justforfun_ ]�U  �]�U  @]�U    ]�U  � ]�U  �b�,�  �9&/       Birthday     �\�U  ��\�U  @�\Some_stuffs_Some_stuffs_ �U  @�\�U  ��\�U  p�\�U  �\�U  �e�,�  �:&/       Appointment P�[�U  п[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��[�U  99h�,�  s;&/       Birthday                       Some_stuffs_Some_stuffs_                                     D m�,�  �<&/      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             
���,�  u_&/       Some_stuffs �7]�U   8]�U  �8]This_stuffs_This_stuffs_ �U   ;]�U  �;]�U  �<]�U   =]�U  ���,�  �d&/       Some_stuffs �*[�U  p+[�U  0,[This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  p0[�U  <e
�,�  �d&/      Appointment �+Z�U  �,Z�U  �5ZSome_stuffs_Some_stuffs_ �U  0/Z�U  �/Z�U  �0Z�U  p1Z�U  1z�,�  >e&/       Workout     `[�U   [�U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `[�U  �G��,�  ��&/       Appointment  �]�U  ��]�U   �]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��]�U  @��,�  ��&/       Some_stuffs ��Y�U  ��Y�U  p�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  ����,�  ��&/       Birthday    `�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   �Z�U  ={��,�  ��&/      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �`$�,�  '�&/      Appointment                    Some_stuffs_Some_stuffs_                                     j�0�,�  Q�&/       Meeting     н[�U  ��[�U  P�[justforfun_justforfun_ [�U  ��[�U  P�[�U  ��[�U  P�[�U  �o5�,�  ��&/       Birthday     �Y�U  �Y�U  0�YSome_stuffs_Some_stuffs_ �U  ��Y�U  ��Y�U  P�Y�U  �Y�U  �T��,�  O�&/       Meeting     ��Z�U  ��Z�U  @�ZSome_stuffs_Some_stuffs_ �U   �Z�U  ��Z�U  ��Z�U   �Z�U  �jǱ,�  ��&/       Birthday    �nZ�U  �oZ�U  ppZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �tZ�U  � Ա,�  %�&/       Appointment ��Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_ �U   �Z�U  ��Z�U  `�Z�U   �Z�U  ��a�,�  k�&/       Birthday    ��^�U  ��^�U  @�^Some_stuffs_Some_stuffs_ �U  ��^�U   �^�U  ��^�U   �^�U   �t�,�  4&/       Some_stuffs @�[�U  ��[�U  ��[justforfun_justforfun_ _ �U  @�[�U  ��[�U  @�[�U  ��[�U  ��,�  �(&/      Birthday     �[�U  ��[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��[�U  *K�,�  	)&/       Workout     �[�U  [�U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  #[�U  �r�,�  a+&/       Some_stuffs                    justforfun_justforfun_                                       J3��,�  ]M&/       Meeting     @{]�U   |]�U  �|]This_stuffs_This_stuffs_ �U  �~]�U  @]�U   �]�U  ��]�U  Xї�,�  �M&/       Meeting ffs 0�X�U  ��X�U  ��Xjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ��X�U  U蝳,�  VO&/      Birthday    ��Z�U  `�Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �Z�U  �p*�,�  Ps&/       Workout     �d^�U  e^�U  �e^justforfun_justforfun_ ^�U  �g^�U  @h^�U  �h^�U  @i^�U  H+>�,�  ]x&/       Workout     p�\�U  �\�U  p�\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��\�U  4Է�,�  ��&/      Appointment 0TY�U   VY�U  @YYSome_stuffs_Some_stuffs_ �U  paY�U  0bY�U  �eY�U  `fY�U  yXǴ,�  {�&/       Birthday fs  eZ�U  �eZ�U  �fZThis_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  pkZ�U  "1ɴ,�  ��&/       Birthday    @Z]�U  �Z]�U  `[]Some_stuffs_Some_stuffs_ �U  �]]�U  `^]�U  �^]�U  `_]�U  �UV�,�  �&/       Appointment ��\�U  @�\�U  ��\justforfun_justforfun_ _ �U  p�\�U  �\�U  ��\�U   �\�U  �}_�,�  n�&/       Workout     �\�U  ��\�U  p�\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�\�U  d�h�,�  ��&/      Workout ent ��Z�U  p�Z�U  0�ZSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  ��Z�U  ʢm�,�  �&/       Workout ffs  �\�U  ��\�U  @�\Some_stuffs_Some_stuffs_ �U  @�\�U   �\�U  ��\�U  ��\�U  �	�,�  ��&/       Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ���,�  e�&/       Workout     @SZ�U   TZ�U  �TZSome_stuffs_Some_stuffs_ �U  �WZ�U  @XZ�U   YZ�U  �YZ�U  6*��,�  B�&/      Birthday    �P\�U  PQ\�U  �Q\justforfun_justforfun_ \�U  PT\�U  �T\�U  PU\�U  �U\�U  +߄�,�  �&/       Appointment �[�U  `[�U   [This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �[�U  ���,�  &/      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ғ��,�  �&/       Workout     �[�U  �[�U   [Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p8[�U  iE��,�  �&/       Appointment p�Y�U  0�Y�U  0�YSome_stuffs_Some_stuffs_ �U   �Y�U  ��Y�U  ��Y�U  p�Y�U  �%�,�  �6&/      Workout  U  ��^�U  @�^�U  ��^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��^�U  ��,�  �\&/      Birthday    0 ]�U  � ]�U  0]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p]�U  �r��,�  �]&/       Some_stuffs �eY�U  `fY�U  �iYThis_stuffs_This_stuffs_ �U  �sY�U  `tY�U  xY�U  �xY�U  qǷ,�  `&/       Birthday    ��\�U   �\�U  ��\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @�\�U  ��O�,�  �&/       Meeting     �E[�U  0F[�U  �F[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �K[�U  JS�,�  �&/       Some_stuffs `^�U  �^�U  `^This_stuffs_This_stuffs_ �U  `^�U   ^�U  �^�U   ^�U  4~Z�,�  &/      Some_stuffs �|Y�U  P}Y�U   �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  QDn�,�  Ҋ&/       Workout      �Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�Z�U  ����,�  ~�&/      Some_stuffs ��[�U  0�[�U  ��[Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  0�[�U  �惹,�  ��&/      Some_stuffs �y\�U  �z\�U   {\justforfun_justforfun_ \�U  @}\�U  �}\�U  @~\�U  �~\�U  ���,�  �&/       Workout     �Z�U  @Z�U  PZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  PZ�U   &��,�  �&/       Workout �U  0�Y�U  �Y�U  ��YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  �	��,�  �&/       Birthday    �[�U  ��[�U  �[justforfun_justforfun_ [�U  ��[�U  �[�U  ��[�U  ��[�U  �!�,�  Y�&/      Workout     �Y�U  `Y�U  �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �&Y�U  q7�,�  ��&/       Workout     �1Y�U  �2Y�U  5Yjustforfun_justforfun_ Y�U  �;Y�U  `<Y�U  @?Y�U  AY�U  �Y��,�  � &/      Birthday    �\�U  ��\�U  �\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��\�U  h;˺,�  �%&/       Appointment  �Y�U  ��Y�U  ��Yjustforfun_justforfun_ Z�U  �Z�U  `Z�U   Z�U  �Z�U  X�O�,�  �G&/       Appointment @�[�U  ��[�U  @�[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��[�U  Х�,�  �n&/       Birthday U   �Z�U  �Z�U  `�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Z�U  Y�,�  �o&/       Appointment 0�Z�U  � [�U  `�ZSome_stuffs_Some_stuffs_ �U  ��Z�U  `�Z�U   �Z�U  ��Z�U  ����,�  o�&/       Meeting ffs ��\�U  0�\�U  ��\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P�\�U  Lֆ�,�  A�&/      Appointment 0�X�U  ��X�U  ��Xjustforfun_justforfun_ X�U  ��X�U  ��X�U  ��X�U  ��X�U  �U��,�  �&/       Birthday    0�]�U  ��]�U  p�]Some_stuffs_Some_stuffs_ �U  �]�U  p�]�U  �]�U  p�]�U  
��,�  �&/       Appointment �V^�U   W^�U  �W^Some_stuffs_Some_stuffs_ �U  �Y^�U  pZ^�U  �Z^�U  p[^�U  ሚ�,�  L�&/       Birthday    0TY�U   VY�U  @YYThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  `fY�U  ���,�  g�&/      Meeting     �Y�U  `Y�U  �YSome_stuffs_Some_stuffs_ �U  �"Y�U  `#Y�U  �%Y�U  �&Y�U  ���,�  d�&/      Appointment ��[�U  @�[�U  ��[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �[�U  ɖ��,�  ��&/       Workout     0�[�U  ��[�U  ��[Some_stuffs_Some_stuffs_ �U  0�[�U  Ь[�U  0�[�U  �[�U  �5�,�  n&/       Appointment [�U  �[�U  �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  [�U  ʿ?�,�  -
&/       Meeting �U  �}]�U  @~]�U  �~]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��]�U  � F�,�  �&/      Birthday nt �O\�U  PP\�U  �P\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �T\�U  ���,�  �/&/      Appointment p�Z�U  0�Z�U   �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  ��b�,�  �T&/       Workout                        justforfun_justforfun_                                       !Vd�,�  U&/       Appointment �0Z�U  p1Z�U  02ZSome_stuffs_Some_stuffs_ �U  �4Z�U  0?Z�U  7Z�U  �7Z�U  ~!t�,�  Y&/      Workout  U  p	]�U  0
]�U  �
]justforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U  �]�U  b��,�  �{&/       Meeting     pP[�U  0Q[�U  �Q[Some_stuffs_Some_stuffs_ �U  pT[�U  �T[�U  �U[�U  0V[�U  ��,�  ��&/      Meeting     02Z�U  �2Z�U  p3ZThis_stuffs_This_stuffs_ �U  7Z�U  �7Z�U  P8Z�U  9Z�U  ��,�  ?�&/       Appointment ��\�U  @�\�U   �\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��\�U  m9��,�  u�&/      Meeting     @�[�U  ��[�U  ��[This_stuffs_This_stuffs_ �U   �[�U  ��[�U  ��[�U   �[�U  躩�,�  a�&/       Some_stuffs ��Z�U  ��Z�U  0�Zjustforfun_justforfun_ Z�U  `�Z�U   �Z�U  ��Z�U  `�Z�U  IE7�,�  ��&/       Workout     �^�U  ��^�U  �^justforfun_justforfun_ ^�U  P�^�U  г^�U  ��^�U  �^�U  <�F�,�  ��&/      Birthday    @�Z�U  ��Z�U  ��ZSome_stuffs_Some_stuffs_ �U  ��Z�U   �Z�U   �Z�U  ��Z�U  $���,�  ��&/      Some_stuffs p�Y�U  0�Y�U  0�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�Y�U  ���,�  ��&/       Appointment �Z�U  �Z�U  PZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Z�U  ���,�  N�&/       Some_stuffs  �Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�Z�U  ��Y�,�  � &/      Some_stuffs  �]�U  ��]�U   �]This_stuffs_This_stuffs_ �U   �]�U  ��]�U  ��]�U  `�]�U  �,b�,�  " &/       Meeting     `�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_ �U  `[�U   [�U  �[�U  `[�U  2��,�  �> &/       Birthday     %_�U  �%_�U  0&_This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  *_�U  �z��,�  a@ &/       Birthday    `�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �Z�U  ��,�  �C &/      Appointment ��Z�U  ��Z�U  p�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �Z�U  ���,�  j &/       Birthday    �Q[�U  pR[�U  0S[Some_stuffs_Some_stuffs_ �U  �U[�U  0V[�U  �V[�U  �W[�U  �Ϟ�,�  1j &/      Appointment @q\�U   r\�U  �r\This_stuffs_This_stuffs_ �U  @u\�U   v\�U  �v\�U   w\�U  �&�,�  Ќ &/       Meeting �U  ppZ�U  0qZ�U  p}ZThis_stuffs_This_stuffs_ �U  0tZ�U  �tZ�U  puZ�U  0vZ�U  }F;�,�  ?� &/      Workout     ��Z�U   �Z�U   �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `�Z�U  !h��,�  T� &/       Some_stuffs 0�[�U  �[�U  p�[justforfun_justforfun_ [�U  0�[�U  ��[�U  0�[�U  ��[�U  kJ��,�  � &/       Appointment ��^�U   �^�U  ��^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `�^�U  "U��,�  t� &/       Appointment `�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_ �U  `�Z�U  ��Z�U  `�Z�U   �Z�U  D���,�  ̻ &/      Birthday    p�Z�U  0�Z�U  ��ZSome_stuffs_Some_stuffs_ �U  ��Z�U  ��Z�U  p�Z�U  ��Z�U  ��c�,�  /� &/       Birthday fs `�\�U  ��\�U  ��\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��\�U  ��p�,�  �� &/       Workout     �Z�U  �Z�U  �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Z�U  ,�s�,�  M� &/      Birthday U   YZ�U  �YZ�U  �ZZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �_Z�U  ����,�  � !&/       Birthday    @VZ�U   WZ�U  �WZThis_stuffs_This_stuffs_ �U  �ZZ�U  @[Z�U   \Z�U  pgZ�U  ���,�  a!&/       Meeting                        Some_stuffs_Some_stuffs_                                     ����,�  !&/      Meeting                        Some_stuffs_Some_stuffs_                                     Z��,�  '!&/       Birthday U  ��Z�U  p�Z�U  0�ZSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ��Z�U  !���,�  �(!&/       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             R���,�  �*!&/       Birthday    �C]�U  D]�U  �D]justforfun_justforfun_ ]�U  �F]�U  0G]�U  �G]�U  0H]�U  x[��,�  [+!&/       Birthday    �[�U  `[�U   [This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �[�U  �
-�,�  6S!&/       Birthday     �[�U  ��[�U  @�[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��[�U  �x��,�  )w!&/      Birthday    xY�U  �xY�U  �|Yjustforfun_justforfun_ Y�U  ��Y�U  ��Y�U  p�Y�U  0�Y�U  4�M�,�  "�!&/      Appointment                    This_stuffs_This_stuffs_                                     Dc��,�  ��!&/      Birthday                       This_stuffs_This_stuffs_                                     ���,�  7�!&/       Workout     �fZ�U  0rZ�U  �gZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �lZ�U  ���,�  �"&/       Birthday    �KZ�U  pLZ�U  0MZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ]Z�U  �.��,�  d9"&/       Meeting     �[\�U  P\\�U   ]\justforfun_justforfun_ \�U  @�\�U  ��\�U  �`\�U  0a\�U  ����,�  (?"&/      Some_stuffs  �Y�U  �Y�U  0�YThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  �Y�U  �q��,�  �?"&/       Birthday    �$Z�U  p-Z�U  &Zjustforfun_justforfun_ Z�U  )Z�U  �)Z�U  P*Z�U  +Z�U  ���,�  �?"&/       Appointment `�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  �K�,�  @a"&/       Birthday    �Z�U  `�Z�U  �ZThis_stuffs_This_stuffs_ �U  `�Z�U   �Z�U  оZ�U  P�Z�U  �L�,�  �a"&/       Birthday    �L[�U  pM[�U  �8[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p=[�U  �Gj�,�  i"&/      Meeting      Z�U  �Z�U  �Zjustforfun_justforfun_ Z�U  �Z�U  �Z�U  �Z�U  pZ�U  W��,�  �"&/      Birthday    �BZ�U  PCZ�U  DZSome_stuffs_Some_stuffs_ �U  GZ�U  �GZ�U  �QZ�U  �RZ�U  � �,�  ��"&/       Meeting                        This_stuffs_This_stuffs_                                     ���,�  {�"&/      Some_stuffs P^\�U  �^\�U  @�\This_stuffs_This_stuffs_ �U  �a\�U  �b\�U  pc\�U  �c\�U  �� �,�  9�"&/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             y�$�,�  [�"&/       Birthday    DZ�U  �DZ�U  �EZSome_stuffs_Some_stuffs_ �U  �QZ�U  �RZ�U  �HZ�U  �IZ�U  �$&�,�  ��"&/      Meeting     [�U  �[�U  P[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P[�U  �|W�,�  �(#&/      Meeting                        This_stuffs_This_stuffs_                                     Q�e�,�  r,#&/       Birthday U  ppZ�U  0qZ�U  p}ZSome_stuffs_Some_stuffs_ �U  0tZ�U  �tZ�U  puZ�U  0vZ�U  ���,�  �S#&/      Some_stuffs                    Some_stuffs_Some_stuffs_                                     �c�#-�  0�-&/      Appointment ��X�U  ��X�U  0�XSome_stuffs_Some_stuffs_ �U   �X�U  ��X�U  ��X�U  @�X�U  ���#-�  ��-&/       Workout     P�Y�U  �Y�U  ��YSome_stuffs_Some_stuffs_ �U   �Y�U  ��Y�U  ��Y�U  ��Y�U  ���#-�  z�-&/       Meeting     pX[�U  0Y[�U  �Y[This_stuffs_This_stuffs_ �U  0\[�U  �\[�U  �][�U  p^[�U  0�>$-�  ~$.&/       Meeting ffs �3[�U  p4[�U  �4[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  pM[�U  �J$-�  �'.&/       Meeting     �`\�U  0a\�U  �a\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �e\�U  �YK$-�  �'.&/      Workout     �m]�U  @n]�U   o]Some_stuffs_Some_stuffs_ �U  @q]�U  �q]�U  @r]�U  �r]�U  B_L$-�  (.&/       Some_stuffs �Z�U  ��Z�U  p�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  =��$-�  �H.&/      Birthday    �Z�U  @Z�U    ZThis_stuffs_This_stuffs_ �U   #Z�U  �#Z�U  �$Z�U  p-Z�U  z�$-�  �M.&/       Workout ffs P�\�U  Н\�U  ��\justforfun_justforfun_ _ �U  �\�U  ��\�U   �\�U  ��\�U  `p�$-�  �O.&/       Birthday U  �e[�U   f[�U  �f[justforfun_justforfun_ [�U  @i[�U  �i[�U  @j[�U  �j[�U  �^%-�  Nn.&/      Appointment ��Y�U  ��Y�U  �Yjustforfun_justforfun_ Y�U  0�Y�U  �Y�U  ��Y�U  @�Y�U  �l%-�  �q.&/       Some_stuffs ��Z�U  `�Z�U   �Zjustforfun_justforfun_ Z�U  `�Z�U   �Z�U  ��Z�U  ��Z�U  �&�%-�  ��.&/       Birthday    �BZ�U  PCZ�U  DZjustforfun_justforfun_ Z�U  GZ�U  �GZ�U  �QZ�U  �RZ�U  �1&-�  k�.&/       Some_stuffs �A[�U  0B[�U  �B[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �G[�U  J&-�  ��.&/       Meeting     0TY�U   VY�U  @YYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `fY�U  |2&-�  ��.&/      Meeting �U   �Y�U  ��Y�U  ��Yjustforfun_justforfun_ Y�U  P�Y�U  �Y�U  ��Y�U  ��Y�U  ��&-�  �.&/      Birthday    �Z�U  �Z�U  `ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �%Z�U  ���&-�  y�.&/       Some_stuffs �G\�U  PH\�U  �H\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �L\�U  �&-�  U�.&/       Workout     P�[�U  �[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P�[�U  9�.'-�  �.&/       Birthday                       Some_stuffs_Some_stuffs_                                     \e;'-�  K�.&/      Workout                        This_stuffs_This_stuffs_                                     �'-�  �/&/      Workout     P�Y�U  �Y�U  ��YSome_stuffs_Some_stuffs_ �U   �Y�U  ��Y�U  ��Y�U  ��Y�U  ���'-�  �/&/       Workout     `�Y�U   �Y�U   �YSome_stuffs_Some_stuffs_ �U  p�Y�U  0�Y�U  ��Y�U  ��Y�U  �9`(-�  B3/&/       Some_stuffs 0_[�U  �_[�U  p`[This_stuffs_This_stuffs_ �U  Pz[�U  �z[�U  @d[�U  �d[�U  �W{(-�  3:/&/      Birthday    ��Z�U  p�Z�U  0�ZThis_stuffs_This_stuffs_ �U  p�Z�U  0�Z�U  ��Z�U  0�Z�U  ��(-�  ?Z/&/       Birthday    `�]�U  ��]�U  `�]Some_stuffs_Some_stuffs_ �U  ��]�U   �]�U  ��]�U   �]�U  ��)-�  �_/&/       Some_stuffs  �Y�U  ��Y�U  ��YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `�Y�U  R�)-�  �/&/       Appointment ��Y�U  @�Y�U  ��YSome_stuffs_Some_stuffs_ �U  ��Y�U  `�Y�U    Z�U  � Z�U  �ޛ)-�  �/&/       Some_stuffs ��\�U  @�\�U  ��\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��\�U  $i�)-�  ��/&/      Meeting �U   #Z�U  �#Z�U  �$Zjustforfun_justforfun_ Z�U  �'Z�U  P(Z�U  )Z�U  �)Z�U  9�)-�  ��/&/       Some_stuffs 0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��X�U  ��1*-�  z�/&/       Meeting     �D]�U  E]�U  �E]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `I]�U  �zB*-�  ��/&/       Some_stuffs �Z�U  ��Z�U  0�Zjustforfun_justforfun_ Z�U  �Z�U  ��Z�U  @�Z�U  ��Z�U  X��*-�  ��/&/       Appointment EY�U  �EY�U  �HYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   VY�U  ��*-�  ��/&/      Appointment 0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  �?\+-�  ��/&/       Birthday    �Y�U  `Y�U  �YThis_stuffs_This_stuffs_ �U  �"Y�U  `#Y�U  �%Y�U  �&Y�U  c!c+-�  ��/&/       Birthday    ��[�U  P�[�U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��[�U  Q�j+-�  ��/&/       Appointment ��[�U  P�[�U  �[This_stuffs_This_stuffs_ �U  ��[�U  `�[�U  �\�U  P\�U  ��w+-�  ��/&/      Birthday    EY�U  �EY�U  �HYThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   VY�U  ���+-�  �0&/       Meeting     ��]�U  @�]�U  ��]This_stuffs_This_stuffs_ �U  ��]�U  ��]�U  �]�U  ��]�U  <0,-�  �!0&/      Some_stuffs [�U  �[�U  �[Some_stuffs_Some_stuffs_ �U  P[�U  [�U  �[�U  [�U  �V�,-�  �F0&/      Appointment �cZ�U  `dZ�U   eZThis_stuffs_This_stuffs_ �U  �gZ�U  phZ�U  0iZ�U  �iZ�U   '<--�  �q0&/       Workout     0�Z�U  ��Z�U  0�ZSome_stuffs_Some_stuffs_ �U  ��Z�U  0�Z�U  �Z�U  ��Z�U  X}�--�  G�0&/       Appointment 0�X�U  ��X�U  ��Xjustforfun_justforfun_ X�U  ��X�U  ��X�U  ��X�U  ��X�U  ��--�  ��0&/      Birthday    ��Z�U  ��Z�U  `�Zjustforfun_justforfun_ Z�U   �Z�U  ��Z�U   �Z�U  ��Z�U  2��--�  >�0&/       Some_stuffs                    justforfun_justforfun_                                       ̊b.-�  �0&/      Workout     5Y�U  �5Y�U  P8YSome_stuffs_Some_stuffs_ �U  @?Y�U  AY�U  EY�U  �EY�U  ��.-�  ��0&/      Appointment @u^�U  �u^�U  @v^This_stuffs_This_stuffs_ �U  �x^�U  `y^�U  �y^�U  `z^�U  �M/-�  E�0&/       Meeting �U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��X�U  �N�/-�  �1&/      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_              ڗ/-�  @1&/       Birthday    �&[�U  0'[�U  �'[justforfun_justforfun_ [�U  �*[�U  p+[�U  0,[�U  �,[�U  � �0-�  �V1&/      Appointment 0TY�U   VY�U  @YYThis_stuffs_This_stuffs_ �U  paY�U  0bY�U  �eY�U  `fY�U  ��0-�  vX1&/       Appointment �_�U  `_�U  �_This_stuffs_This_stuffs_ �U  �_�U  `_�U  �_�U  `_�U  ��P1-�  }1&/       Some_stuffs PU\�U  �U\�U  PV\justforfun_justforfun_ \�U  Y\�U  �Y\�U  PZ\�U  [\�U  <�a1-�  w�1&/      Meeting                        justforfun_justforfun_                                       �>i1-�  d�1&/       Some_stuffs pP[�U  0Q[�U  �Q[This_stuffs_This_stuffs_ �U  pT[�U  �T[�U  �U[�U  0V[�U  �On1-�  ��1&/       Workout     `�]�U  ��]�U  `�]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �]�U  -�1-�  $�1&/      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �E�1-�  �1&/       Birthday nt `�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `[�U  j�2-�  q�1&/       Appointment `_^�U  ��^�U  ``^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  d^�U  }�2-�  ?�1&/      Appointment �KZ�U  pLZ�U  0MZThis_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U   ]Z�U  &�2-�  ��1&/       Workout �U  0TY�U   VY�U  @YYSome_stuffs_Some_stuffs_ �U  paY�U  0bY�U  �eY�U  `fY�U  ��2-�  ��1&/       Meeting     @s]�U  �s]�U  @t]This_stuffs_This_stuffs_ �U  �v]�U  �w]�U   x]�U  �x]�U  8d3-�  ��1&/      Some_stuffs 0�X�U  ��X�U  ��Xjustforfun_justforfun_ X�U  ��X�U  ��X�U  ��X�U  ��X�U  �,3-�  ��1&/       Workout �U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  �f3-�  ��1&/       Meeting �U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��X�U  PT$3-�  ��1&/       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ��)3-�  E�1&/       Workout                        This_stuffs_This_stuffs_                                     c303-�  ��1&/       Workout     �%Y�U  �&Y�U  )Yjustforfun_justforfun_ Y�U  �1Y�U  �2Y�U  5Y�U  �5Y�U  �13-�  ?�1&/       Birthday    PAZ�U  �AZ�U  �BZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �GZ�U  �|63-�  x�1&/       Some_stuffs `\�U   \�U  �\Some_stuffs_Some_stuffs_ �U  0\�U  �\�U  �\�U  p\�U  �]�3-�  A2&/       Birthday                       justforfun_justforfun_                                       ���3-�  �2&/      Some_stuffs  �Y�U  ��Y�U  ��YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Z�U  2u�3-�   2&/       Birthday    @(]�U  �(]�U  p)]Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   -]�U   �H4-�  �?2&/       Birthday    ��X�U  @�X�U   YSome_stuffs_Some_stuffs_ �U  PY�U  Y�U   	Y�U  �	Y�U  �]L4-�  �@2&/      Appointment ��Y�U  ��Y�U  �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @�Y�U  �ZS4-�  eB2&/       Appointment �Y�U  `Y�U  �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �&Y�U  3�g4-�  �G2&/       Some_stuffs �q[�U  Pr[�U  s[justforfun_justforfun_ [�U  Pu[�U  �u[�U  Pv[�U  w[�U  p��4-�  &g2&/       Some_stuffs P]Y�U  ^Y�U  paYThis_stuffs_This_stuffs_ �U  �iY�U  �jY�U  @oY�U   pY�U  ��4-�  *g2&/       Birthday    p�Z�U  ��Z�U  ��ZSome_stuffs_Some_stuffs_ �U  p�Z�U  �Z�U  ��Z�U  p�Z�U  ��4-�  zi2&/      Birthday     ]\�U  �]\�U  P^\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �b\�U  ��4-�  �l2&/       Appointment ``^�U  a^�U  �a^Some_stuffs_Some_stuffs_ �U  �c^�U  d^�U  �d^�U  e^�U  �<_-�  �>=&/       Some_stuffs ��[�U  p�[�U  �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �[�U  �K_-�  �B=&/      Birthday U    Z�U  � Z�U  �!ZThis_stuffs_This_stuffs_ �U  �$Z�U  p-Z�U  &Z�U  �&Z�U   w�_-�  �c=&/       Birthday    p�[�U  �[�U  P�[justforfun_justforfun_ [�U  ��[�U  P�[�U  �[�U  б[�U  ���_-�  He=&/      Meeting     ��\�U   �\�U  ��\Some_stuffs_Some_stuffs_ �U  P�\�U  Щ\�U  p�\�U  0�\�U  j5�_-�  �e=&/       Birthday nt ��]�U  `�]�U   �]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��]�U  �=o`-�  �=&/      Appointment ��\�U  @�\�U  ��\This_stuffs_This_stuffs_ �U  ��\�U  p�\�U  0�\�U  ��\�U  ��a-�  e�=&/       Meeting     ��[�U  ��[�U  @�[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @�[�U  �a-�  ��=&/      Appointment �yZ�U  0zZ�U  �zZSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  ��Z�U  }��a-�  ?�=&/      Some_stuffs  �Z�U  ��Z�U   �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  �G�a-�  ��=&/       Some_stuffs  �\�U  ��\�U   �\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �\�U  ��a-�  ��=&/       Meeting     5Y�U  �5Y�U  P8YThis_stuffs_This_stuffs_ �U  @?Y�U  AY�U  EY�U  �EY�U  �'9b-�  X>&/       Workout      \�U  �\�U  `\Some_stuffs_Some_stuffs_ �U   \�U  �\�U  `\�U   \�U  �:b-�  �>&/       Meeting     �<Z�U  P=Z�U  >Zjustforfun_justforfun_ Z�U  PAZ�U  �AZ�U  �BZ�U  PCZ�U  f�@b-�  @>&/      Birthday      ]�U  � ]�U  0!]This_stuffs_This_stuffs_ �U  0#]�U  �#]�U  �Q]�U  pR]�U  p��b-�  �+>&/       Birthday nt �]�U  0]�U  �]This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  0]�U  8R|c-�  U>&/       Workout     �\�U  ��\�U  @�\Some_stuffs_Some_stuffs_ �U  ��\�U   �\�U  ��\�U  @�\�U  "yd-�  �x>&/       Workout     ��]�U  p�]�U  ��]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��]�U  y�d-�  �y>&/       Workout ffs �][�U  p^[�U  0_[justforfun_justforfun_ [�U  �a[�U  0b[�U  Pz[�U  �z[�U  p d-�  �{>&/       Workout     `�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_ �U  ��Z�U  ��Z�U  @�Z�U   �Z�U  �Ѡd-�  ��>&/      Meeting �U  0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��X�U  "Ţd-�  t�>&/       Workout     �,\�U  P-\�U  .\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �2\�U  	�d-�  �>&/       Birthday U  �4[�U  p5[�U  �5[justforfun_justforfun_ [�U  �L[�U  pM[�U  �8[�U  p9[�U  1-*e-�  �>&/       Workout  fs PV\�U  W\�U  �W\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P\\�U  @�0e-�  ��>&/       Appointment ��]�U   �]�U  ��]justforfun_justforfun_ ]�U   �]�U  ��]�U   �]�U  ��]�U  ��e-�  ��>&/       Workout     �!Z�U  @"Z�U   #ZThis_stuffs_This_stuffs_ �U  &Z�U  �&Z�U  �'Z�U  P(Z�U  ��^f-�  -?&/       Some_stuffs PU\�U  �U\�U  PV\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  [\�U  1<`f-�  ~?&/       Some_stuffs 0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��X�U  3�af-�  �?&/       Some_stuffs EY�U  �EY�U  �HYjustforfun_justforfun_ Y�U  �PY�U  @QY�U  0TY�U   VY�U  H�df-�  �?&/       Appointment �Y�U  `Y�U  �YThis_stuffs_This_stuffs_ �U  �"Y�U  `#Y�U  �%Y�U  �&Y�U  �!�f-�  �7?&/       Meeting     p�Z�U  ��Z�U  ��ZSome_stuffs_Some_stuffs_ �U  p�Z�U  �Z�U  ��Z�U  p�Z�U  `-�f-�  8?&/       Birthday     YZ�U  �YZ�U  �ZZSome_stuffs_Some_stuffs_ �U  �]Z�U  `^Z�U   _Z�U  �_Z�U  ��g-�  ??&/      Meeting     t[�U  �t[�U  Pu[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �y[�U  BI�g-�  H^?&/       Meeting     ��\�U  `�\�U   �\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `�\�U  ��g-�  �a?&/      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �5�g-�  ne?&/       Meeting      �[�U  ��[�U  @�[justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ��[�U  ~�3h-�  �?&/      Workout      �\�U  ��\�U  ��\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0�\�U  ��3h-�  +�?&/       Workout     0JZ�U  �JZ�U  �KZSome_stuffs_Some_stuffs_ �U  pNZ�U  0OZ�U  �OZ�U  �PZ�U  ��3h-�  +�?&/       Appointment ��Z�U  0�Z�U  �ZSome_stuffs_Some_stuffs_ �U  ��Z�U  p�Z�U  0�Z�U  ��Z�U  %��h-�  ��?&/      Some_stuffs @s]�U  �s]�U  @t]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �x]�U  l�h-�  U�?&/       Workout     0,[�U  �,[�U  p-[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �1[�U  ��_i-�  ��?&/      Appointment 0TY�U   VY�U  @YYSome_stuffs_Some_stuffs_ �U  paY�U  0bY�U  �eY�U  `fY�U  Rqgi-�  ��?&/       Some_stuffs @_�U  �_�U  p_Some_stuffs_Some_stuffs_ �U  �	_�U  `
_�U  �
_�U  `_�U  3�mi-�  ��?&/       Birthday    `�]�U   �]�U  ��]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��]�U  �1oi-�  ��?&/       Some_stuffs 0]�U  �]�U  p]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p]�U  q��i-�  ��?&/       Workout     xY�U  �xY�U  �|YSome_stuffs_Some_stuffs_ �U  ��Y�U  ��Y�U  p�Y�U  0�Y�U  J�j-�  }@&/       Some_stuffs �~Z�U  0Z�U  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0�Z�U  ,hj-�  -@&/      Meeting     �Z�U  @Z�U  PZThis_stuffs_This_stuffs_ �U  PZ�U  �Z�U  �Z�U  PZ�U  �ٟj-�  �(@&/       Some_stuffs @r]�U  �r]�U  @s]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �w]�U  �ˤj-�  0*@&/       Workout     0\�U  �\�U  �\This_stuffs_This_stuffs_ �U  �\�U  0\�U  �\�U  p\�U  D9"k-�  LJ@&/      Birthday    ��X�U  @�X�U   YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �	Y�U  �,�k-�  �o@&/      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �_�k-�  r@&/       Meeting  U   B^�U  �B^�U   C^justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  G^�U  q�k-�  Fv@&/       Appointment ��X�U  ��X�U  0�XSome_stuffs_Some_stuffs_ �U   �X�U  ��X�U  ��X�U  @�X�U  �pl-�  @&/       Appointment &Z�U  �&Z�U  �'ZSome_stuffs_Some_stuffs_ �U  P*Z�U  +Z�U  �+Z�U  �,Z�U  @C�l-�  ��@&/       Birthday    ��Y�U  ��Y�U  `�Yjustforfun_justforfun_ Y�U  ��Y�U  ��Y�U  p�Y�U  0�Y�U  �l-�  9�@&/      Birthday    ��[�U  @�[�U  ��[This_stuffs_This_stuffs_ �U  @�[�U  ��[�U  ��[�U  @�[�U  ��m-�  ��@&/      Some_stuffs  �Z�U  ��Z�U   �ZThis_stuffs_This_stuffs_ �U  ��Z�U  `�Z�U  ��Z�U  ��Z�U  A��m-�  �@&/       Appointment �,]�U   -]�U  �-]justforfun_justforfun_ ]�U  0]�U  �0]�U  1]�U  �1]�U  y%n-�  �A&/       Meeting �U  0�X�U  ��X�U  ��Xjustforfun_justforfun_ X�U  ��X�U  ��X�U  ��X�U  ��X�U  01n-�  �A&/       Workout     p�Z�U  0�Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  x�n-�  �5A&/       Appointment                    This_stuffs_This_stuffs_                                     �@�n-�  �5A&/      Birthday fs pe\�U  �e\�U  pf\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �j\�U  b�Io-�  �ZA&/       Appointment @�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Z�U  �
Ko-�  �ZA&/       Meeting     DZ�U  �DZ�U  �EZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �IZ�U  ��Ro-�  �\A&/       Workout �U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  ��do-�  �aA&/      Workout     P*\�U  +\�U  �+\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P0\�U  �;�o-�  ځA&/       Birthday U  �QZ�U  �RZ�U  �HZSome_stuffs_Some_stuffs_ �U  �KZ�U  pLZ�U  0MZ�U  �MZ�U  ���o-�  ��A&/       Appointment  �]�U  ��]�U   �]justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ��]�U  ���o-�  Z�A&/       Appointment `�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_ �U  ��Z�U  `�Z�U   �Z�U  ��Z�U  :l p-�  S�A&/       Meeting     0�Z�U  ��Z�U  `�ZThis_stuffs_This_stuffs_ �U  @�Z�U   �Z�U  ��Z�U  ��Z�U  `*yp-�  <�A&/       Birthday                       justforfun_justforfun_                                       ��p-�  ��A&/      Meeting      �Y�U  ��Y�U  ��YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Z�U  )�p-�  �A&/       Some_stuffs p�Y�U  0�Y�U  0�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p�Y�U  ���p-�  C�A&/       Some_stuffs 0�[�U  Ь[�U  0�[justforfun_justforfun_ [�U  �[�U  ��[�U  0�[�U  �[�U  �q-�  ��A&/      Birthday    xY�U  �xY�U  �|YThis_stuffs_This_stuffs_ �U  ��Y�U  ��Y�U  p�Y�U  0�Y�U  �'q-�  ��A&/       Some_stuffs 0]�U  �]�U  p	]justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  �]�U  YQ˚-�  �}L&/       Workout     �%Y�U  �&Y�U  )YSome_stuffs_Some_stuffs_ �U  �1Y�U  �2Y�U  5Y�U  �5Y�U  �W՚-�  X�L&/       Workout     Л\�U  ��\�U  P�\justforfun_justforfun_ \�U  ��\�U  `�\�U  �\�U  ��\�U  �'�-�  /�L&/      Meeting     �jZ�U  pkZ�U  0lZSome_stuffs_Some_stuffs_ �U  �nZ�U  �oZ�U  ppZ�U  0qZ�U  ��{�-�  ��L&/       Appointment ��^�U  `�^�U  �^This_stuffs_This_stuffs_ �U  �^�U  ��^�U  @�^�U  ��^�U  D��-�  ��L&/      Appointment ��Y�U  ��Y�U  �YSome_stuffs_Some_stuffs_ �U  `�Y�U   �Y�U  ��Y�U  `�Y�U  ���-�  ��L&/       Workout  U  0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ��X�U  X�	�-�  G�L&/       Birthday                       This_stuffs_This_stuffs_                                     �$�-�  ��L&/      Birthday    p_�U   _�U  �_justforfun_justforfun_ _�U  �
_�U  `_�U  �_�U  `_�U  X/��-�  ��L&/       Meeting �U    Z�U  � Z�U  �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Z�U  �.��-�  �L&/      Workout     @2]�U  �2]�U  `3]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   7]�U  �/�-�  eM&/       Meeting     ppZ�U  0qZ�U  p}ZSome_stuffs_Some_stuffs_ �U  0tZ�U  �tZ�U  puZ�U  0vZ�U  �VA�-�  M&/      Meeting ffs ��Y�U  p�Y�U  ��YSome_stuffs_Some_stuffs_ �U  �Y�U  ��Y�U   �Y�U  �Y�U  �J�-�  N!M&/       Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             c+P�-�  �"M&/       Appointment 0�[�U  ��[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0�[�U  ��˝-�  �BM&/       Workout �U  �Z�U  ��Z�U  p�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �Z�U  "�-�  @IM&/       Some_stuffs �Z�U  @Z�U  PZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  PZ�U  z�-�  {IM&/       Meeting     �<^�U  P=^�U  �=^This_stuffs_This_stuffs_ �U   @^�U  �@^�U   A^�U  �A^�U  ��g�-�  ejM&/       Meeting �U  �U[�U  0V[�U  �V[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �[[�U  1�m�-�  �kM&/       Appointment p�\�U  0�\�U  ��\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �\�U  o�-�  NlM&/      Appointment  �^�U  ��^�U   �^Some_stuffs_Some_stuffs_ �U   �^�U  ��^�U   �^�U  ��^�U  �;~�-�  0pM&/       Some_stuffs  C^�U  �C^�U  `D^This_stuffs_This_stuffs_ �U  �F^�U  G^�U  �G^�U  H^�U  ��-�  d�M&/      Appointment �+Z�U  �,Z�U  �5ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p1Z�U  aK�-�  ܖM&/       Workout     `[�U   [�U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `[�U  P��-�  �M&/       Meeting      �Y�U  ��Y�U  ��YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  \�)�-�  ��M&/      Meeting �U  p�Y�U  0�Y�U  0�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�Y�U  �q/�-�  �M&/       Birthday nt 0]�U  �]�U  p]This_stuffs_This_stuffs_ �U  �]�U  0]�U  �]�U  p]�U  ��@�-�  ��M&/       Some_stuffs 0�[�U  ��[�U  0�[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��[�U  �XǠ-�  �N&/       Appointment `\�U   \�U  �\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p\�U  D�Π-�  �N&/      Birthday                       Some_stuffs_Some_stuffs_                                     rp�-�  D1N&/      Birthday    @d[�U  �d[�U  �e[This_stuffs_This_stuffs_ �U   h[�U  �h[�U  @i[�U  �i[�U  )�-�  IVN&/       Some_stuffs  �[�U  ��[�U  @�[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��[�U  ,"�-�  m[N&/      Appointment �Z�U  ��Z�U  p�ZSome_stuffs_Some_stuffs_ �U  0�Z�U  ��Z�U  @�Z�U   �Z�U  �鐢-�  {N&/      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             @MC�-�  ȨN&/       Some_stuffs �1Y�U  �2Y�U  5YThis_stuffs_This_stuffs_ �U  �;Y�U  `<Y�U  @?Y�U  AY�U   "£-�  @�N&/       Workout ent ��Y�U  p�Y�U  ��YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Y�U  <e�-�  ��N&/      Some_stuffs  �]�U  ��]�U   �]This_stuffs_This_stuffs_ �U  `�]�U  ��]�U  `�]�U   �]�U  �_�-�  �O&/      Meeting      _Z�U  �_Z�U  �`ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �eZ�U  ���-�  �=O&/       Birthday nt  	Y�U  �	Y�U  �YSome_stuffs_Some_stuffs_ �U  �Y�U  `Y�U  �Y�U  `Y�U  ����-�  c@O&/       Appointment ��Y�U  ��Y�U  �YSome_stuffs_Some_stuffs_ �U  `�Y�U   �Y�U  ��Y�U  `�Y�U  = ��-�  �CO&/      Appointment pe\�U  �e\�U  pf\This_stuffs_This_stuffs_ �U  �h\�U  �i\�U   j\�U  �j\�U  �#�-�  _eO&/       Appointment 0�[�U  �[�U  p�[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��[�U  t=5�-�  �iO&/      Workout     0MZ�U  �MZ�U  pNZSome_stuffs_Some_stuffs_ �U  �\Z�U   ]Z�U  @SZ�U   TZ�U   �˦-�  `�O&/       Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             S7ͦ-�  ��O&/       Some_stuffs 0\�U  �\�U  0\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @>\�U  )Oئ-�  ��O&/       Birthday U   �Z�U  ��Z�U   �ZThis_stuffs_This_stuffs_ �U  ��Z�U  `�Z�U  ��Z�U  ��Z�U  ��٦-�  �O&/      Appointment ��]�U  p�]�U  ��]Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ��]�U  I�V�-�  ݳO&/       Workout     p�Z�U  0�Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0�Z�U  R0`�-�  R�O&/       Some_stuffs  [�U  �[�U  `[Some_stuffs_Some_stuffs_ �U   [�U  �[�U  `	[�U   
[�U  ��p�-�  ��O&/      Some_stuffs �Z�U  ��Z�U   �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Z�U  �-�  ��O&/      Workout     ��Z�U  ��Z�U  @�ZThis_stuffs_This_stuffs_ �U  `�Z�U   �Z�U  ��Z�U  `�Z�U  �0�-�  ��O&/       Appointment ��Z�U  0�Z�U  �ZThis_stuffs_This_stuffs_ �U  �Z�U  p�Z�U  ��Z�U  ��Z�U  <q��-�  wP&/      Workout ffs @�[�U  ��[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �[�U  ��*�-�  �+P&/       Some_stuffs �'[�U  p([�U  0)[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �-[�U  a�/�-�  �,P&/       Appointment  bZ�U  �bZ�U  �cZSome_stuffs_Some_stuffs_ �U  �fZ�U  0rZ�U  �gZ�U  phZ�U  jK:�-�  �/P&/       Appointment P�\�U  Щ\�U  p�\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��\�U  ©-�  uRP&/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��ө-�  �VP&/       Some_stuffs @�]�U  ��]�U  @�]justforfun_justforfun_ ]�U  ��]�U  @�]�U  ��]�U  @�]�U  �qK�-�  �uP&/      Workout     P�]�U  ��]�U  ��]This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  ��]�U  �n[�-�  �yP&/       Some_stuffs ��Z�U  `�Z�U   �ZThis_stuffs_This_stuffs_ �U  ��Z�U  `�Z�U  ��Z�U  ` [�U  ^�-�  _zP&/       Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             L�-�  �P&/      Appointment ��Z�U  ��Z�U  p�Zjustforfun_justforfun_ Z�U  0�Z�U  ��Z�U  `�Z�U   �Z�U  A+�-�  ��P&/       Workout     �?Z�U  �@Z�U  PAZThis_stuffs_This_stuffs_ �U  DZ�U  �DZ�U  �EZ�U  PFZ�U  "$��-�  ԡP&/       Some_stuffs `[]�U   \]�U  �\]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ``]�U  mD��-�  U�P&/      Appointment p"\�U  �"\�U  �#\Some_stuffs_Some_stuffs_ �U  &\�U  �&\�U  P'\�U  (\�U  b֛�-�  ��P&/       Workout ent  �Y�U  ��Y�U  ��YThis_stuffs_This_stuffs_ �U  ��Y�U  ��Y�U  �Y�U  ��Y�U  ���-�  �P&/       Workout     �Y�U  `Y�U  �Yjustforfun_justforfun_ Y�U  �"Y�U  `#Y�U  �%Y�U  �&Y�U  ���-�  k�P&/       Workout ffs �[�U  �[�U  `[justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  �$[�U  ���-�  ~�P&/      Meeting �U  �zZ�U  �{Z�U  p|ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0�Z�U  �k�-�  j�[&/       Appointment 0�Z�U  ��Z�U  p�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Z�U  �$x�-�  ��[&/       Workout     p|Z�U  �|Z�U  �~ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  �|�-�  ��[&/      Some_stuffs �rZ�U  psZ�U  0tZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �xZ�U  ���-�  x�[&/       Some_stuffs  	Y�U  �	Y�U  �YThis_stuffs_This_stuffs_ �U  �Y�U  `Y�U  �Y�U  `Y�U  в��-�  ��[&/       Meeting     �|Y�U  P}Y�U   �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  �y�-�  ��[&/      Meeting     P*Z�U  +Z�U  �+Zjustforfun_justforfun_ Z�U  �-Z�U  �.Z�U  0/Z�U  �/Z�U  侞�-�  \&/      Meeting �U   �Y�U  ��Y�U  ��YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Z�U  �/�-�  95\&/      Meeting �U  PT\�U  �T\�U  PU\This_stuffs_This_stuffs_ �U  �W\�U  PX\�U  Y\�U  �Y\�U  (|��-�  �a\&/       Some_stuffs P4\�U  �4\�U  P5\This_stuffs_This_stuffs_ �U  �7\�U  P8\�U  �8\�U  �9\�U  ��i�-�  ��\&/       Birthday    �%Y�U  �&Y�U  )YThis_stuffs_This_stuffs_ �U  �1Y�U  �2Y�U  5Y�U  �5Y�U  $Em�-�  x�\&/      Some_stuffs �0Z�U  p1Z�U  02ZSome_stuffs_Some_stuffs_ �U  �4Z�U  0?Z�U  7Z�U  �7Z�U  ����-�  �\&/       Birthday     Z�U  �Z�U  �Zjustforfun_justforfun_ Z�U  �Z�U  �Z�U  �Z�U  pZ�U  ��-�   �\&/       Meeting     �Z�U  pZ�U  0	ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @Z�U  Bc�-�  ��\&/       Meeting ffs ��\�U  p$]�U  ��\justforfun_justforfun_ _ �U  �\�U  ��\�U  �\�U  ��\�U  �*�-�  >�\&/      Workout �U  ��X�U  @�X�U   Yjustforfun_justforfun_ Y�U  PY�U  Y�U   	Y�U  �	Y�U  h���-�  �\&/       Workout ent ��]�U  P�]�U  И]This_stuffs_This_stuffs_ �U  К]�U  P�]�U  Л]�U  ��]�U  �׫�-�  �\&/      Meeting     ��Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  j9�-�  D�\&/      Birthday    p�[�U  0�[�U  �[This_stuffs_This_stuffs_ �U  p�[�U  �[�U  ��[�U  p�[�U  *A�-�  @�\&/       Workout     ��[�U  �[�U  ��[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��[�U  ��K�-�  � ]&/       Some_stuffs �QZ�U  �RZ�U  �HZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �MZ�U  ���-�  , ]&/       Birthday    �sY�U  `tY�U  xYSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ��Y�U  L3��-�  a#]&/      Birthday    �BZ�U  PCZ�U  DZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �RZ�U  ipd�-�  �H]&/       Appointment �&[�U  0'[�U  �'[Some_stuffs_Some_stuffs_ �U  �*[�U  p+[�U  0,[�U  �,[�U  x�s�-�  �L]&/       Birthday    0�Z�U  ��Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p�Z�U  ����-�  n]&/      Birthday    ��]�U  ��]�U   �]Some_stuffs_Some_stuffs_ �U   �]�U  ��]�U   �]�U  ��]�U  �q �-�  �p]&/       Birthday fs  �]�U  ��]�U   �]This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U   �]�U  ꥞�-�  A�]&/       Some_stuffs @VZ�U   WZ�U  �WZjustforfun_justforfun_ _ �U  �ZZ�U  @[Z�U   \Z�U  pgZ�U  ���-�  ��]&/      Birthday    г[�U  ��[�U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �[�U  1.��-�  ��]&/       Workout ffs  A]�U  �A]�U  `B]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  F]�U  K%�-�  ��]&/      Meeting     �%Y�U  �&Y�U  )YThis_stuffs_This_stuffs_ �U  �1Y�U  �2Y�U  5Y�U  �5Y�U  ɻ4�-�  ��]&/       Some_stuffs ��^�U   �^�U  ��^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `�^�U  $��-�  �]&/      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             )(��-�  )�]&/       Appointment ��[�U  p�[�U  �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �[�U  �V�-�  �	^&/       Birthday    ��]�U  @�]�U  ��]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��]�U  1i�-�  �^&/       Birthday                       justforfun_justforfun_ _                                     ��v�-�  ^&/      Workout �U  0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  ���-�  s2^&/      Some_stuffs  �Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�Z�U  P���-�  �W^&/       Birthday    ��Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Z�U  �%�-�  B�^&/       Birthday U  @(]�U  �(]�U  p)]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   -]�U  <T%�-�  W�^&/      Some_stuffs �F[�U  �G[�U  pH[Some_stuffs_Some_stuffs_ �U  0K[�U  �K[�U  c[�U  �c[�U  Q�=�-�  ��^&/       Appointment  �\�U  ��\�U  ��\This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  0�\�U  Ec��-�  ��^&/      Meeting �U  0TY�U   VY�U  @YYSome_stuffs_Some_stuffs_ �U  paY�U  0bY�U  �eY�U  `fY�U   ��-�  �^&/       Some_stuffs 0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  �S�-�  ��^&/       Some_stuffs P�[�U  �[�U  н[justforfun_justforfun_ [�U  ��[�U  �[�U  ��[�U  P�[�U  �HS�-�  ��^&/       Birthday nt ��Z�U  0�Z�U  ��Zjustforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U   �Z�U  �Bn�-�  ��^&/       Appointment �[�U  P[�U  [Some_stuffs_Some_stuffs_ �U  �[�U  �[�U  [�U  �[�U  ��r�-�  ��^&/       Meeting �U  �%Y�U  �&Y�U  )YThis_stuffs_This_stuffs_ �U  �1Y�U  �2Y�U  5Y�U  �5Y�U  ,#t�-�  �^&/      Birthday                       Some_stuffs_Some_stuffs_                                     ���-�  �^&/       Workout      �Y�U  ��Y�U  ��YThis_stuffs_This_stuffs_ �U  0�Y�U  ��Y�U   �Y�U  ЕY�U  (��-�  ��^&/       Some_stuffs ��Y�U  ��Y�U  �YSome_stuffs_Some_stuffs_ �U  `�Y�U   �Y�U  ��Y�U  `�Y�U  $���-�  �_&/      Workout                        Some_stuffs_Some_stuffs_                                     z��-�  �_&/       Birthday     �Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_ �U  ��Z�U  `�Z�U   �Z�U  �Z�U  �J��-�  a"_&/       Birthday    �Y�U  `Y�U  �YSome_stuffs_Some_stuffs_ �U  �"Y�U  `#Y�U  �%Y�U  �&Y�U  U)�-�  �E_&/      Appointment ��X�U  ��X�U  0�Xjustforfun_justforfun_ X�U   �X�U  ��X�U  ��X�U  @�X�U  ���-�  Xi_&/       Birthday     _Z�U  �_Z�U  �`ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �eZ�U  ዾ�-�  ,l_&/       Workout     ��Y�U  ��Y�U  �YThis_stuffs_This_stuffs_ �U  `�Y�U   �Y�U  ��Y�U  `�Y�U  N��-�  !p_&/      Birthday    @k[�U  �k[�U  �l[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   q[�U  �Mf�-�  �_&/      Meeting     0MZ�U  �MZ�U  pNZThis_stuffs_This_stuffs_ �U  �\Z�U   ]Z�U  @SZ�U   TZ�U  �u��-�  p�_&/       Meeting ent p�^�U  ��^�U  p�^This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U   �^�U  l���-�  չ_&/      Workout     �Z�U  ��Z�U  p�Zjustforfun_justforfun_ Z�U  0�Z�U  ��Z�U  @�Z�U   �Z�U  z�-�  �_&/      Some_stuffs                    justforfun_justforfun_                                       A��-�  ��_&/       Workout     p�Z�U  �Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  C�"�-�  �`&/       Some_stuffs ��\�U  `�\�U  ��\justforfun_justforfun_ \�U   �\�U  ��\�U   �\�U  ��\�U  A�+�-�  (`&/       Birthday    0�\�U  ��\�U  0 ]This_stuffs_This_stuffs_ �U  p]�U  0]�U  �]�U  0]�U  �/�-�  	`&/      Birthday    �Z�U  @Z�U  PZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  PZ�U  ��2�-�  `&/       Birthday    ��[�U  P�[�U  �[Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  �[�U  �}��-�  A0`&/       Workout     �Z�U  �Z�U  PZThis_stuffs_This_stuffs_ �U  Z�U  �Z�U  �Z�U  �Z�U  ����-�  g1`&/      Birthday                       justforfun_justforfun_                                       �I�-�  =T`&/      Appointment �[�U  [�U  �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  #[�U  0SS�-�  �V`&/       Workout                        justforfun_justforfun_                                       ��.�  Zk&/      Meeting     �A[�U  0B[�U  �B[Some_stuffs_Some_stuffs_ �U  �E[�U  0F[�U  �F[�U  �G[�U  ��.�  �,k&/      Meeting ffs �$]�U  p%]�U  �%]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �)]�U  (�.�  �1k&/       Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             dj1.�  <Pk&/       Birthday nt @2]�U  �2]�U  `3]justforfun_justforfun_ _ �U  `5]�U  �5]�U  �6]�U   7]�U  V�4.�  Qk&/      Birthday U  ��[�U  P�[�U  г[This_stuffs_This_stuffs_ �U  P�[�U  ж[�U  P�[�U  з[�U  �k6.�  �Qk&/       Meeting     0TY�U   VY�U  @YYSome_stuffs_Some_stuffs_ �U  paY�U  0bY�U  �eY�U  `fY�U  s�I.�  �Vk&/       Some_stuffs �o\�U  �p\�U  @q\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   v\�U  �mQ.�  nXk&/       Workout     ��Y�U  ��Y�U  p�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  ��.�  �wk&/       Appointment �\Z�U   ]Z�U  @SZjustforfun_justforfun_ Z�U  @VZ�U   WZ�U  �WZ�U  @XZ�U  �K�.�  �yk&/       Some_stuffs 0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��X�U  P�v.�  ��k&/       Some_stuffs ��[�U  p�[�U  0�[justforfun_justforfun_ [�U  0�[�U  ��[�U  p�[�U  0�[�U  �y.�  D�k&/      Meeting     ��]�U  `�]�U   �]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �]�U  �C.�  ��k&/       Birthday    ��Z�U  `�Z�U   �Zjustforfun_justforfun_ Z�U  ��Z�U  ��Z�U  0�Z�U  ��Z�U  M=.�  ��k&/      Some_stuffs P�[�U  п[�U  ��[Some_stuffs_Some_stuffs_ �U  ��[�U  P�[�U  �[�U  ��[�U  ��.�  ��k&/       Workout     ��^�U  �^�U  ��^justforfun_justforfun_ ^�U  ��^�U  @�^�U  ��^�U  @�^�U  !c�.�  4�k&/       Meeting     ��\�U   �\�U  ��\Some_stuffs_Some_stuffs_ �U  p�\�U  ��\�U  ��\�U  @�\�U  p�.�  ��k&/      Appointment �Z�U  @Z�U  PZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  PZ�U  P�C.�  �l&/       Birthday    ��X�U  @�X�U   YThis_stuffs_This_stuffs_ �U  PY�U  Y�U   	Y�U  �	Y�U  �jF.�  8l&/       Birthday     �Z�U  ��Z�U  `�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   [�U  ��L.�  �l&/      Birthday nt �*[�U  p+[�U  0,[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p0[�U  ��.�  �:l&/       Meeting     0�[�U  Ь[�U  0�[justforfun_justforfun_ [�U  �[�U  ��[�U  0�[�U  �[�U  ��.�  �=l&/       Workout     ��\�U  p�\�U  �\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �\�U  �/�.�  �Bl&/      Appointment �d]�U  0e]�U  �e]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �i]�U  �0g.�  %dl&/       Appointment  �]�U  ��]�U  `�]Some_stuffs_Some_stuffs_ �U  ��]�U   �]�U  ��]�U   �]�U  \�k.�  Kel&/      Workout �U  0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��X�U  �Wt.�  �gl&/       Meeting     �Z�U  ��Z�U   �Zjustforfun_justforfun_ _ �U  оZ�U  P�Z�U  0�Z�U  �Z�U  ��.�  �jl&/       Some_stuffs �=[�U  �>[�U  p?[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  pC[�U  ��.�  �jl&/       Meeting     `\�U  �\�U  `\justforfun_justforfun_ \�U  �\�U  `\�U   \�U  �\�U  ��.�  Z�l&/      Some_stuffs @�\�U  ��\�U  p�\This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  Н\�U  ��.�  o�l&/       Workout                        This_stuffs_This_stuffs_                                     �Ǯ.�  �l&/       Birthday    �x\�U  @y\�U  �y\justforfun_justforfun_ _ �U   |\�U  �|\�U  @}\�U  �}\�U  ,X0.�  -�l&/      Some_stuffs �&[�U  0'[�U  �'[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �,[�U  �=5.�  n�l&/       Birthday fs P�^�U  ��^�U  P�^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `�^�U  ��B.�  ��l&/       Appointment �+]�U   ,]�U  �,]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �0]�U  Q��.�  ��l&/       Workout      \�U  �\�U  `\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �\�U  t��.�  jm&/      Appointment ��Y�U  `�Y�U   �YThis_stuffs_This_stuffs_ �U  p�Y�U  0�Y�U  ��Y�U  ��Y�U  T�f.�  �(m&/      Meeting     �Q[�U  pR[�U  0S[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �W[�U  �r.�  �+m&/       Workout     �g^�U  @h^�U  �h^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �l^�U  �_�.�  -Nm&/       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ���.�  �Om&/      Meeting     ��Y�U  ��Y�U  �YSome_stuffs_Some_stuffs_ �U  `�Y�U   �Y�U  ��Y�U  `�Y�U  �q.�  �Pm&/       Some_stuffs                    Some_stuffs_Some_stuffs_                                     �^�.�  tm&/       Some_stuffs ��Z�U  ��Z�U  `�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `�Z�U  ��".�  P�m&/       Meeting     �\�U  p\�U  0\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �\�U  @ $.�  ��m&/       Appointment  �Y�U  ��Y�U  ��YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  1L+.�  ~�m&/       Meeting     0�Z�U  ��Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p�Z�U  �?.�  ��m&/      Workout �U  �>_�U  @?_�U  �?_justforfun_justforfun_ _�U  �A_�U  pB_�U  �B_�U  pC_�U  )��.�  I�m&/       Workout     ppZ�U  0qZ�U  p}ZSome_stuffs_Some_stuffs_ �U  0tZ�U  �tZ�U  puZ�U  0vZ�U  $��.�  X�m&/      Some_stuffs                    Some_stuffs_Some_stuffs_                                     Q,a.�  ��m&/       Workout      �Y�U  ��Y�U  ��Yjustforfun_justforfun_ Z�U  �Z�U  `Z�U   Z�U  �Z�U  ފl.�  ��m&/      Birthday    �6\�U  7\�U  �7\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P<\�U  Ёr.�  B�m&/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �r�.�  �n&/      Appointment ��Z�U  ��Z�U  0�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0�Z�U  8��.�  Sn&/       Birthday    �g\�U  0h\�U  �h\Some_stuffs_Some_stuffs_ �U  @k\�U  �k\�U  @l\�U  �l\�U  ��.�  �6n&/      Birthday nt 0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��X�U  �a�.�  k8n&/       Appointment 0JZ�U  �JZ�U  �KZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �PZ�U  ��.�  p<n&/       Workout     ��Z�U  p�Z�U  0�ZSome_stuffs_Some_stuffs_ �U  p�Z�U  0�Z�U  ��Z�U  0�Z�U  � .�  :^n&/      Meeting                        This_stuffs_This_stuffs_                                     1�4.�  ~cn&/       Meeting       Z�U  � Z�U  �!ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �&Z�U  X�.�  �n&/       Birthday    �Y�U  `Y�U  �YSome_stuffs_Some_stuffs_ �U  �"Y�U  `#Y�U  �%Y�U  �&Y�U  ��.�  s�n&/      Some_stuffs �\�U  ��\�U  @�\justforfun_justforfun_ _ �U  ��\�U   �\�U  ��\�U  @�\�U  Z��.�  ��n&/       Workout ffs �jZ�U  pkZ�U  0lZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0qZ�U  ��.�  �n&/       Workout     �Z�U  PZ�U  ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Z�U  ô�.�  x�n&/       Some_stuffs   \�U  � \�U  `\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   \�U  hzk .�  �n&/       Meeting �U  0MZ�U  �MZ�U  pNZjustforfun_justforfun_ Z�U  �\Z�U   ]Z�U  @SZ�U   TZ�U  7�� .�  ~�n&/       Birthday fs ��Z�U  `�Z�U   �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Z�U  TB� .�  ��n&/       Birthday    �[�U  �[�U  P[justforfun_justforfun_ _ �U  �[�U  �[�U   [�U  � [�U  :.� .�  ��n&/       Appointment  Z�U  �Z�U  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pZ�U  �Z� .�  ��n&/      Appointment �]Z�U  `^Z�U   _ZThis_stuffs_This_stuffs_ �U   bZ�U  �bZ�U  �cZ�U  `dZ�U  c�!.�  |�n&/       Workout     L]�U  �L]�U  M]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �P]�U  ��!.�  ��n&/       Meeting     ��Y�U  ��Y�U   �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  UA!.�  ��n&/       Meeting     ��\�U  @�\�U  ��\justforfun_justforfun_ \�U  ��\�U  @�\�U  ��\�U  ��\�U  ��!.�  Z�n&/       Appointment ��]�U  P�]�U  И]Some_stuffs_Some_stuffs_ �U  К]�U  P�]�U  Л]�U  ��]�U  �N�!.�  ��n&/       Workout     �!Z�U  @"Z�U   #ZSome_stuffs_Some_stuffs_ �U  &Z�U  �&Z�U  �'Z�U  P(Z�U  �!.�  5�n&/       Appointment ��\�U  �\�U  ��\This_stuffs_This_stuffs_ �U  ��\�U  `�\�U  ��\�U  `�\�U  �:�!.�   o&/       Birthday    ��X�U  ��X�U  0�XThis_stuffs_This_stuffs_ �U   �X�U  ��X�U  ��X�U  @�X�U  ���!.�  so&/      Some_stuffs `	[�U   
[�U  �
[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `[�U  �Y$".�  �#o&/       Meeting ffs  Z�U  �Z�U  �ZSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  pZ�U  ��0".�  'o&/       Birthday    `�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_ �U  ��Z�U  p�Z�U  0�Z�U  ��Z�U  I"�".�  �Ho&/       Appointment  �\�U  �\�U  ��\This_stuffs_This_stuffs_ �U  ��\�U  @�\�U  P�\�U  Щ\�U  N��".�  aIo&/      Workout ffs 9^�U  �9^�U  p:^justforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U  P>^�U  ���".�  �Ko&/       Workout ffs  �\�U  �\�U  ��\justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  Щ\�U  mI#.�  �no&/       Appointment `	[�U   
[�U  �
[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `[�U  %Z#.�  8so&/      Birthday    �[�U  P[�U  [Some_stuffs_Some_stuffs_ �U  �[�U  �[�U  [�U  �[�U  5b�#.�  B�o&/      Meeting     0JZ�U  �JZ�U  �KZjustforfun_justforfun_ Z�U  pNZ�U  0OZ�U  �OZ�U  �PZ�U   ��#.�  ��o&/       Meeting     �"[�U  #[�U  �#[Some_stuffs_Some_stuffs_ �U  �&[�U  0'[�U  �'[�U  p([�U  I�M.�  �Ez&/       Some_stuffs �U[�U  0V[�U  �V[This_stuffs_This_stuffs_ �U  �Y[�U  pZ[�U  0[[�U  �[[�U  l¡M.�  Fz&/      Appointment xY�U  �xY�U  �|YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0�Y�U  b/�M.�  \Mz&/       Appointment  �]�U  ��]�U   �]Some_stuffs_Some_stuffs_ �U  ��]�U  `�]�U  ��]�U  `�]�U  ���N.�  :�z&/       Some_stuffs 0�]�U  �]�U  p�]This_stuffs_This_stuffs_ �U  p�]�U  �]�U  p�]�U  �]�U  ��N.�  ��z&/      Some_stuffs PN\�U  �N\�U  �O\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �S\�U  |�uO.�  ߽z&/      Appointment puZ�U  0vZ�U  �vZSome_stuffs_Some_stuffs_ �U  �yZ�U  0zZ�U  �zZ�U  �{Z�U  R�uO.�  �z&/       Meeting     EY�U  �EY�U  �HYjustforfun_justforfun_ Y�U  �PY�U  @QY�U  0TY�U   VY�U  �G�O.�  Z�z&/       Workout     �Z�U  ��Z�U  @�ZThis_stuffs_This_stuffs_ �U  ��Z�U  ��Z�U  p�Z�U  ��Z�U  t��P.�  j
{&/      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             r��P.�  �{&/       Meeting ent @�\�U  ��\�U  �`\This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  �d\�U  )��P.�  	{&/       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �)9Q.�  s1{&/      Birthday    ��Z�U  0�Z�U  �ZThis_stuffs_This_stuffs_ �U  �Z�U  p�Z�U  ��Z�U  ��Z�U  !&OQ.�  7{&/       Birthday    @�\�U  ��\�U  ��\justforfun_justforfun_ \�U  ��\�U  @�\�U  ��\�U  @�\�U  �8�Q.�  y\{&/       Meeting     p`[�U  �`[�U  �a[Some_stuffs_Some_stuffs_ �U  @d[�U  �d[�U  �e[�U   f[�U  ���Q.�  /^{&/      Workout                        This_stuffs_This_stuffs_                                     aR.�  5}{&/       Meeting                        This_stuffs_This_stuffs_                                     �FlR.�  �{&/      Meeting ffs `[�U  �[�U  �[justforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U  P[�U  �NuR.�  b�{&/       Some_stuffs t[�U  �t[�U  Pu[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �y[�U  ��R.�  �{&/       Workout     ��[�U  p�[�U  0�[This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  ��[�U  �l�R.�  |�{&/      Workout ffs �[�U  ��[�U  ��[justforfun_justforfun_ _ �U  �[�U  ��[�U  P�[�U  ��[�U  F S.�  ��{&/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �S.�  է{&/       Workout     V]�U  �V]�U  PW]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   \]�U  I�S.�  ��{&/       Meeting     0tZ�U  �tZ�U  puZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0zZ�U  �`S.�  !�{&/       Workout     ��Z�U  ��Z�U  @�ZThis_stuffs_This_stuffs_ �U   �Z�U  ��Z�U  ��Z�U   �Z�U  �S.�  6�{&/       Meeting      �Y�U  ��Y�U  ��YSome_stuffs_Some_stuffs_ �U  P�Y�U  �Y�U  ��Y�U  ��Y�U  ly�S.�  u�{&/      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �6T.�  G�{&/      Workout     �I[�U  pJ[�U  0K[Some_stuffs_Some_stuffs_ �U  N[�U  �N[�U  pO[�U  �O[�U  ���T.�  �|&/       Meeting     �}]�U  @~]�U  �~]justforfun_justforfun_ ]�U  0�]�U  ��]�U  0�]�U  ��]�U  �%�T.�  n|&/       Birthday    ��\�U  ��\�U  @�\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �\�U  ���T.�  �|&/       Birthday nt ��Z�U  `�Z�U  ��ZSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  �[�U  ���T.�  ~ |&/      Meeting                        justforfun_justforfun_                                       tI�U.�  Ji|&/      Birthday      Z�U  � Z�U  �!ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �&Z�U  �B�U.�  j|&/       Birthday    0�[�U  ��[�U  ��[This_stuffs_This_stuffs_ �U  0�[�U  ��[�U  ��[�U  0�[�U  P��V.�  ��|&/       Birthday    [�U  �[�U  P[This_stuffs_This_stuffs_ �U  [�U  �[�U  �[�U  P[�U  Ai�V.�  H�|&/       Appointment �Y�U  `Y�U  �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �&Y�U  �ťV.�  �|&/      Meeting     �B\�U  @C\�U   D\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  PH\�U  ���V.�  d�|&/       Meeting     ��Z�U  p�Z�U  0�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �Z�U  T�3W.�  V�|&/      Appointment                    justforfun_justforfun_                                       D�W.�  l�|&/      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             y"�W.�  ��|&/       Birthday     h[�U  �h[�U  @i[This_stuffs_This_stuffs_ �U  @k[�U  �k[�U  �l[�U   m[�U  �hhX.�  L}&/       Meeting     0\�U  �\�U  �\Some_stuffs_Some_stuffs_ �U  �\�U  0\�U  �\�U  p\�U  � mX.�  y	}&/       Birthday    ��Z�U  ��Z�U  @�Zjustforfun_justforfun_ Z�U  @�Z�U   �Z�U  ��Z�U  ��Z�U  �&wX.�  }&/      Some_stuffs p�\�U  ��\�U  ��\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��\�U  |k�X.�  _+}&/      Birthday    �%Y�U  �&Y�U  )YSome_stuffs_Some_stuffs_ �U  �1Y�U  �2Y�U  5Y�U  �5Y�U  �� Y.�  E/}&/       Some_stuffs  �]�U  ��]�U   �]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �]�U  وY.�  #R}&/      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��1Z.�  m}}&/       Meeting     0�Y�U  �Y�U  ��YSome_stuffs_Some_stuffs_ �U  P�Y�U  �Y�U  ��Y�U  ��Y�U  U�BZ.�  ��}&/      Meeting     0K[�U  �K[�U  c[justforfun_justforfun_ [�U  pO[�U  �O[�U  pP[�U  0Q[�U  ���Z.�  N�}&/       Birthday    �5Z�U  P6Z�U  �-ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �2Z�U  AY�Z.�  H�}&/       Meeting     ��[�U  �[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P�[�U  ٓV[.�  W�}&/       Birthday    0TY�U   VY�U  @YYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `fY�U  *QX[.�  ��}&/       Appointment `�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  4�`[.�  ��}&/      Workout �U  0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��X�U  S�k[.�  ��}&/       Workout     0]�U  �]�U  0]justforfun_justforfun_ ]�U  �
]�U  0]�U  �]�U  �]�U  Qx�[.�  R�}&/       Birthday    @�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Z�U  T�	\.�  6�}&/      Workout �U  0�X�U  ��X�U  ��Xjustforfun_justforfun_ X�U  ��X�U  ��X�U  ��X�U  ��X�U  䍋\.�  p~&/      Workout     �+Z�U  �,Z�U  �5ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p1Z�U  �W].�  �<~&/       Meeting     p%[�U  0&[�U  �&[justforfun_justforfun_ _ �U  0)[�U  �)[�U  �*[�U  p+[�U  �*].�  @~&/      Some_stuffs p�Y�U  0�Y�U  0�YSome_stuffs_Some_stuffs_ �U   �Y�U  ��Y�U  ��Y�U  p�Y�U  ,b�].�  mc~&/      Birthday U  ��Y�U  ��Y�U  p�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  &��].�  �c~&/       Some_stuffs �[�U  е[�U  P�[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��[�U  �].�   e~&/       Appointment p\�U  �\�U  �\This_stuffs_This_stuffs_ �U  \�U  �\�U  @ \�U  � \�U  �+�].�  i~&/       Workout �U  p�Z�U  ��Z�U  ��ZThis_stuffs_This_stuffs_ �U  `�Z�U   �Z�U  ��Z�U  ��Z�U  ���].�  k~&/       Some_stuffs ��\�U  @�\�U  ��\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��\�U  Jc�].�  ]k~&/       Birthday    �Y�U  `Y�U  �YSome_stuffs_Some_stuffs_ �U  �"Y�U  `#Y�U  �%Y�U  �&Y�U  ��].�  �k~&/       Meeting     @�[�U  ��[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P�[�U  �h^.�  ��~&/      Workout     �\�U  ��\�U  0�\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �]�U  ���^.�  l�~&/       Appointment p�Y�U  0�Y�U  0�YSome_stuffs_Some_stuffs_ �U   �Y�U  ��Y�U  ��Y�U  p�Y�U  +��^.�  )�~&/       Birthday fs �[�U  �[�U   [This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p8[�U  ��^.�  ��~&/       Birthday nt @u]�U   v]�U  �v]justforfun_justforfun_ _ �U   y]�U  �y]�U  @z]�U  �z]�U   �^.�  Է~&/       Some_stuffs ��[�U  0�[�U  �[justforfun_justforfun_ [�U  ��[�U  0�[�U  �[�U  p�[�U  	>�.�  ���&/       Appointment p^�U  0^�U  �^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �_^�U   .K�.�  ��&/       Meeting     ��\�U  ��\�U  0�\justforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U  @�\�U  8��.�  �&/       Appointment pmZ�U  0nZ�U  �nZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  psZ�U  ��t�.�  D؉&/       Some_stuffs ��[�U  p�[�U  0�[justforfun_justforfun_ _ �U  0�[�U  ��[�U  0�[�U  ��[�U  {�.�  �ى&/       Workout     `�]�U  ��]�U  ��]Some_stuffs_Some_stuffs_ �U  ��]�U  p�]�U  ��]�U  ��]�U  �r|�.�  :ډ&/       Some_stuffs �%Y�U  �&Y�U  )YThis_stuffs_This_stuffs_ �U  �1Y�U  �2Y�U  5Y�U  �5Y�U  ��.�  ۉ&/       Some_stuffs P![�U  "[�U  �"[This_stuffs_This_stuffs_ �U  p%[�U  0&[�U  �&[�U  0'[�U  ���.�  lۉ&/       Birthday U  �X_�U   Y_�U  �Y_This_stuffs_This_stuffs_ �U  �[_�U  P\_�U  �\_�U  P]_�U  :���.�  �݉&/       Meeting ent P5\�U  6\�U  �6\justforfun_justforfun_ \�U  �8\�U  �9\�U  P:\�U  ;\�U  H0�.�  }��&/       Some_stuffs                    justforfun_justforfun_                                       ���.�  	�&/      Appointment ��Y�U  ��Y�U  p�Yjustforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U  �Y�U  H���.�  �)�&/       Birthday     �Z�U  ��Z�U  `�ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �Z�U  �o��.�  Z*�&/       Workout     `�Z�U  ��Z�U  `�ZThis_stuffs_This_stuffs_ �U  `�Z�U   �Z�U  ��Z�U  `�Z�U  F-��.�  �*�&/      Some_stuffs  �Y�U  ��Y�U  ��YThis_stuffs_This_stuffs_ �U  0�Y�U  ��Y�U   �Y�U  ЕY�U  IE;�.�  �L�&/       Appointment `�Y�U   �Y�U  ��YThis_stuffs_This_stuffs_ �U  ��Y�U  ��Y�U  p�Y�U  0�Y�U  \LC�.�  �N�&/      Some_stuffs                    Some_stuffs_Some_stuffs_                                     �"Q�.�  6R�&/       Appointment ��^�U  @�^�U  ��^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��^�U  �o،.�  �t�&/       Some_stuffs                    This_stuffs_This_stuffs_                                     nc�.�  n��&/      Birthday      Z�U  � Z�U  �!ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �&Z�U  �xt�.�  ˜�&/       Meeting     p-[�U  �-[�U  �.[This_stuffs_This_stuffs_ �U  01[�U  �1[�U  �2[�U  03[�U  �t�.�  ~Ŋ&/      Meeting     ��Z�U  ��Z�U  @�ZThis_stuffs_This_stuffs_ �U   �Z�U  ��Z�U  ��Z�U   �Z�U  B|��.�  (�&/       Some_stuffs 0\�U  �\�U  �\justforfun_justforfun_ \�U  �\�U  0\�U  �\�U  p\�U  ݜ��.�  ��&/      Some_stuffs p�Z�U  0�Z�U  ��Zjustforfun_justforfun_ Z�U  0�Z�U  �Z�U  ��Z�U  0�Z�U  �ñ�.�  �&/       Some_stuffs 0�[�U  Ь[�U  0�[Some_stuffs_Some_stuffs_ �U  �[�U  ��[�U  0�[�U  �[�U  �&2�.�  ��&/       Appointment                    This_stuffs_This_stuffs_                                     �?�.�  n�&/      Meeting �U  P�Y�U  �Y�U  ��YSome_stuffs_Some_stuffs_ �U   �Y�U  ��Y�U  ��Y�U  ��Y�U  �bۏ.�  6:�&/       Meeting     �KZ�U  pLZ�U  0MZThis_stuffs_This_stuffs_ �U  �OZ�U  �PZ�U  �\Z�U   ]Z�U  ��ޏ.�  ;�&/       Some_stuffs �1Y�U  �2Y�U  5YThis_stuffs_This_stuffs_ �U  �;Y�U  `<Y�U  @?Y�U  AY�U  9��.�  S=�&/       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             h�r�.�  �`�&/       Some_stuffs N^�U  �N^�U  O^This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  �R^�U  �B~�.�  �c�&/      Workout      �Y�U  �Y�U  0�YSome_stuffs_Some_stuffs_ �U  ��Y�U  ��Y�U  P�Y�U  �Y�U  *���.�  ɂ�&/       Workout     M]�U  �M]�U  PN]This_stuffs_This_stuffs_ �U  PP]�U  �P]�U  PQ]�U  ��]�U  ���.�  g��&/      Meeting     @�[�U   �[�U  ��[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��[�U   ��.�  ���&/       Some_stuffs ��Y�U   �Y�U  ��YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  ɳ��.�  ���&/       Meeting     �sY�U  `tY�U  xYjustforfun_justforfun_ Y�U   �Y�U  ��Y�U  ��Y�U  ��Y�U  �Y��.�  �&/       Meeting  nt �-_�U  ._�U  �._Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  2_�U  _��.�  9��&/      Workout     0�Y�U  ��Y�U  `�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  ��@�.�  G׋&/      Meeting ffs ��[�U  0�[�U  ��[Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ��[�U  �4ǒ.�  ���&/      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             1ns�.�  �%�&/       Workout     �a[�U  0b[�U  Pz[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @g[�U  �kx�.�  '�&/       Some_stuffs ��Y�U  ��Y�U  P�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  (=��.�  It�&/       Appointment `�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  ��!�.�  㓌&/       Meeting �U  ��Y�U  ��Y�U  �YThis_stuffs_This_stuffs_ �U  `�Y�U   �Y�U  ��Y�U  `�Y�U  %�"�.�  8��&/      Some_stuffs  �Y�U  ��Y�U  ��Yjustforfun_justforfun_ Y�U  P�Y�U  �Y�U  ��Y�U  ��Y�U  �'/�.�  V��&/       Appointment ��[�U  �[�U  ��[justforfun_justforfun_ _ his_stuffs_This_stuffs_ �U  ��[�U  )	��.�  ��&/       Meeting ent  �Y�U  ��Y�U  ��YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Z�U  L��.�  �&/      Birthday    @�\�U  �\�U  p�\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �\�U  ���.�  �1�&/       Some_stuffs ��[�U   �[�U  ��[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @�[�U  l���.�  2�&/      Birthday U  �Z�U  �Z�U  PZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Z�U  "z��.�  �3�&/       Appointment ��^�U   �^�U  ��^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0�^�U  9���.�  �8�&/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��*�.�  �Z�&/      Some_stuffs PT\�U  �T\�U  PU\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �Y\�U  �-�.�  �[�&/       Birthday    0\�U  �\�U  p\justforfun_justforfun_ \�U  �\�U  @>\�U  \�U  �\�U  �k<�.�  W_�&/       Appointment ��X�U  P�X�U   �XSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pY�U  �TƘ.�  ���&/       Meeting �U  @SZ�U   TZ�U  �TZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �YZ�U  ��Ș.�  E��&/       Workout     0TY�U   VY�U  @YYjustforfun_justforfun_ Y�U  paY�U  0bY�U  �eY�U  `fY�U  C*Ϙ.�  脍&/       Appointment ��Y�U  ��Y�U   �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  �Ԙ.�  )��&/      Some_stuffs   Z�U  � Z�U  �!ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �&Z�U  ��՘.�  ���&/       Workout ent ��]�U  @�]�U  ��]Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ��]�U  ��V�.�  ���&/       Birthday    0)[�U  �)[�U  �*[justforfun_justforfun_ _ �U  p-[�U  �-[�U  �.[�U  p/[�U  �\�.�  ���&/       Some_stuffs PZ�U  �Z�U  �Zjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U   Z�U  �(c�.�  ˪�&/       Some_stuffs @A\�U   B\�U  �B\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  G\�U  !:f�.�  ���&/       Appointment 0\�U  �\�U  0\Some_stuffs_Some_stuffs_ �U  �\�U  p\�U  �\�U  @>\�U  ���.�  �э&/      Workout ffs �]�U  0]�U  �]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ]�U  ���.�  �Ӎ&/       Appointment `�Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   �Z�U  ʀ�.�  ��&/       Workout     �%Y�U  �&Y�U  )YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �5Y�U  �섚.�  ��&/       Birthday    �\�U  p\�U  0\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �\�U  �c��.�  ���&/       Appointment pNZ�U  0OZ�U  �OZSome_stuffs_Some_stuffs_ �U  @SZ�U   TZ�U  �TZ�U  �UZ�U  @��.�  ���&/       Meeting     ��Z�U  `�Z�U   �Zjustforfun_justforfun_ Z�U  �Z�U  `�Z�U  �Z�U  ��Z�U  G,��.�  (��&/       Meeting     �yZ�U  0zZ�U  �zZjustforfun_justforfun_ Z�U  �~Z�U  0Z�U  �Z�U  ��Z�U  �ᚚ.�  ���&/       Meeting     ��[�U  p�[�U  0�[This_stuffs_This_stuffs_ �U  ��[�U  0�[�U  ��[�U  ��[�U  aP��.�  ���&/       Workout     �Y�U  `Y�U  �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �&Y�U  >���.�  ��&/      Some_stuffs �Y�U  `Y�U  �YThis_stuffs_This_stuffs_ �U  �"Y�U  `#Y�U  �%Y�U  �&Y�U  ��&�.�  p�&/      Birthday    ��X�U  @�X�U   YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �	Y�U  kX��.�  �ɘ&/       Workout     L\�U  �L\�U  PM\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  PQ\�U  y���.�  �͘&/       Appointment �[�U  �[�U  P[justforfun_justforfun_ [�U  �[�U  �[�U   [�U  � [�U  "E��.�  tИ&/       Appointment  �Z�U  ��Z�U  `�Zjustforfun_justforfun_ _ �U  ��Z�U  ��Z�U  `�Z�U   �Z�U  
��.�  �ј&/      Appointment ��X�U  ��X�U  0�XThis_stuffs_This_stuffs_ �U   �X�U  ��X�U  ��X�U  @�X�U  Ī��.�  <��&/      Some_stuffs pmZ�U  0nZ�U  �nZjustforfun_justforfun_ Z�U  p}Z�U  �}Z�U  �rZ�U  psZ�U  d��.�  <�&/       Appointment �]�U  �]�U  `]Some_stuffs_Some_stuffs_ �U  �]�U  @]�U  �]�U  @]�U  *e�.�  I�&/       Meeting     @�[�U  ��[�U  @�[Some_stuffs_Some_stuffs_ �U  ��[�U  @�[�U   �[�U  ��[�U  	��.�  u�&/       Birthday    [�U  �[�U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  [�U  ��.�  x�&/       Workout     �Z�U  ��Z�U  p�ZSome_stuffs_Some_stuffs_ �U  0�Z�U  ��Z�U  @�Z�U   �Z�U  $�!�.�  8�&/      Some_stuffs                    This_stuffs_This_stuffs_                                     ���.�  �B�&/      Appointment _�U  �_�U  _Some_stuffs_Some_stuffs_ �U  p_�U  �_�U  p_�U   _�U  x\��.�  �E�&/       Workout     ��]�U  @�]�U  ��]justforfun_justforfun_ ]�U   �]�U  ��]�U   �]�U  ��]�U  ��5�.�  �e�&/       Birthday    p%[�U  0&[�U  �&[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p+[�U  
�:�.�  g�&/       Meeting     1]�U  �1]�U  @2]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �5]�U  �D�.�  ~i�&/      Appointment �eY�U  `fY�U  �iYSome_stuffs_Some_stuffs_ �U  �sY�U  `tY�U  xY�U  �xY�U  ���.�  ��&/      Birthday                       justforfun_justforfun_                                       ��d�.�  T��&/      Appointment ��Y�U  ��Y�U  P�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Y�U  A��.�  h��&/       Meeting     `�Z�U   �Z�U  ��ZThis_stuffs_This_stuffs_ �U  ��Z�U  `�Z�U   �Z�U  ��Z�U  �L��.�  x��&/       Meeting ffs 0]�U  �]�U  p	]justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  �]�U  �} �.�  Cۙ&/       Appointment  �Y�U  ЕY�U   �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  �$	�.�  zݙ&/      Meeting     �Z�U  pZ�U  0	ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @Z�U  7�.�  ��&/       Some_stuffs ��Z�U  0�Z�U  �ZSome_stuffs_Some_stuffs_ �U  �Z�U  p�Z�U  ��Z�U  ��Z�U  "��.�  ��&/       Meeting                        This_stuffs_This_stuffs_                                     9,��.�  S�&/       Workout     xY�U  �xY�U  �|YSome_stuffs_Some_stuffs_ �U  ��Y�U  ��Y�U  p�Y�U  0�Y�U  2	��.�  ��&/       Meeting     �0^�U  P1^�U  �1^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   6^�U  4H��.�  �&/      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             -�D�.�  M.�&/      Some_stuffs ��[�U  0�[�U  ��[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0�[�U  �bL�.�  :0�&/       Appointment �%Y�U  �&Y�U  )YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �5Y�U  �n��.�  =P�&/      Appointment �<Z�U  P=Z�U  >ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  PCZ�U  /j�.�  dy�&/      Meeting     �QZ�U  �RZ�U  �HZThis_stuffs_This_stuffs_ �U  �KZ�U  pLZ�U  0MZ�U  �MZ�U  ��n�.�  �z�&/       Workout                        This_stuffs_This_stuffs_                                     Pv�.�  |�&/       Birthday    0#]�U  �#]�U  �Q]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �']�U  C�z�.�  �}�&/       Some_stuffs ��[�U  p�[�U  0�[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�[�U  rG|�.�  ~�&/       Birthday    �[�U  ��[�U  P�[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �[�U  ����.�  p��&/      Some_stuffs ��Y�U  ��Y�U  �Yjustforfun_justforfun_ Y�U  `�Y�U   �Y�U  ��Y�U  `�Y�U  � 
�.�  N��&/       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             I՗�.�  �ƚ&/       Birthday    �[�U  �[�U  [Some_stuffs_Some_stuffs_ �U  �[�U  �[�U  P[�U  [�U  |Z��.�  �ƚ&/      Birthday    0TY�U   VY�U  @YYThis_stuffs_This_stuffs_ �U  paY�U  0bY�U  �eY�U  `fY�U  ��E�.�  &�&/      Meeting     �[�U  [�U  �[Some_stuffs_Some_stuffs_ �U  P![�U  "[�U  �"[�U  #[�U  �K�.�  ���&/       Workout     �&^�U  �'^�U   (^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �+^�U  Y;��.�  �&/       Meeting     ��[�U  P�[�U  �[justforfun_justforfun_ [�U  ��[�U  `�[�U   �[�U  ��[�U  *l��.�  ��&/       Meeting     �Z�U  pZ�U  0	ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @Z�U  0���.�  ^�&/       Some_stuffs @�[�U  ��[�U  ��[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��[�U  h�j�.�  1>�&/       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             YEk�.�  G>�&/       Meeting     P8Z�U  9Z�U  �9ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pHZ�U  ���.�  �d�&/       Workout     ��[�U  0�[�U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p�[�U  ��.�  �f�&/       Workout     �4[�U  p5[�U  �5[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p9[�U  �S�.�  h�&/      Workout     �<Z�U  P=Z�U  >ZSome_stuffs_Some_stuffs_ �U  PAZ�U  �AZ�U  �BZ�U  PCZ�U  ����.�  ���&/      Some_stuffs ��Z�U  `�Z�U   �ZSome_stuffs_Some_stuffs_ �U  ��Z�U  ��Z�U  0�Z�U  ��Z�U  Yr��.�  g��&/       Workout     `�Z�U  �Z�U  `�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   �Z�U  z��.�  ۍ�&/       Birthday    ��Y�U  p�Y�U  ��YThis_stuffs_This_stuffs_ �U   �Y�U  �Y�U  0�Y�U  �Y�U  �6�.�  ٳ�&/      Appointment �Z�U  �Z�U  �ZThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  0Z�U  ����.�  0֛&/       Some_stuffs 0JZ�U  �JZ�U  �KZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �PZ�U  ,���.�  �ܛ&/      Workout     �+Z�U  �,Z�U  �5ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p1Z�U  1�V�.�  ���&/       Meeting     ��Z�U   �Z�U  ��ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  �X[�.�  ���&/       Appointment ��\�U  p�\�U  0�\This_stuffs_This_stuffs_ �U  p�\�U  0�\�U  ��\�U  p�\�U  
Qu�.�  u�&/       Some_stuffs `\�U  �\�U  `\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �\�U  �x�.�  '�&/      Workout     �[�U  `[�U   [This_stuffs_This_stuffs_ �U  �[�U  P[�U  [�U  �[�U  p��.�  f%�&/       Meeting                        justforfun_justforfun_                                       ]���.�  �%�&/      Some_stuffs ��\�U  @�\�U  ��\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��\�U  Z���.�  G&�&/       Birthday    ��X�U  ��X�U  0�XThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @�X�U  �O��.�  �'�&/       Appointment ��Z�U  0�Z�U  ��Zjustforfun_justforfun_ [�U  `�Z�U  ��Z�U  `�Z�U   �Z�U  ��.�  �O�&/      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �2 �.�  �r�&/      Some_stuffs M]�U  �M]�U  PN]This_stuffs_This_stuffs_ �U  PP]�U  �P]�U  PQ]�U  ��]�U  x�/�.�  �v�&/       Appointment @z]�U  �z]�U  @{]Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  @]�U  ����.�  h��&/      Appointment �9Z�U  P:Z�U  ;Zjustforfun_justforfun_ Z�U  >Z�U  pHZ�U  �?Z�U  �@Z�U  `��.�  \��&/       Birthday    �zZ�U  �{Z�U  p|ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0�Z�U  ����.�  .��&/       Meeting     0/Z�U  �/Z�U  �0Zjustforfun_justforfun_ Z�U  p3Z�U  04Z�U  �4Z�U  0?Z�U  [���.�  ���&/       Birthday nt p�]�U  �]�U  ��]Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  p�]�U  �9X�.�  �&/      Birthday                       justforfun_justforfun_ _Some_stuffs_Some_stuffs_             qij�.�  Fǜ&/       Birthday U   YZ�U  �YZ�U  �ZZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �_Z�U  Y���.�  ��&/       Some_stuffs �[�U  p�[�U  0�[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �[�U  ���.�  �&/       Appointment  �^�U  ��^�U  P�^justforfun_justforfun_ ^�U  ��^�U   �^�U  ��^�U   �^�U  �d��.�  ��&/       Birthday    �]�U  @]�U  �]Some_stuffs_Some_stuffs_ �U  0!]�U  �!]�U  0"]�U  �"]�U  <�.�  W�&/      Appointment ��Z�U  p�Z�U  0�ZSome_stuffs_Some_stuffs_ �U  ��Z�U  0�Z�U  �Z�U  ��Z�U  �V��.�  �&/       Meeting     ��Z�U  0�Z�U  �Zjustforfun_justforfun_ _ �U  ��Z�U  p�Z�U  0�Z�U  ��Z�U  �՗�.�  p�&/      Meeting     ��Z�U  p�Z�U  0�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Z�U  Q��.�  ��&/       Some_stuffs  �Y�U  ��Y�U  ��YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0�Y�U  S;/�.�  2;�&/       Some_stuffs ��^�U   �^�U  ��^This_stuffs_This_stuffs_ �U  �^�U  `�^�U  �^�U  ��^�U  ��1�.�  �;�&/      Appointment p�Y�U  0�Y�U  0�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�Y�U  ��2�.�  <�&/       Some_stuffs xY�U  �xY�U  �|Yjustforfun_justforfun_ Y�U  ��Y�U  ��Y�U  p�Y�U  0�Y�U  ��6�.�  =�&/       Workout     ��[�U  0�[�U  �[Some_stuffs_Some_stuffs_ �U  ��[�U  0�[�U  �[�U  p�[�U  b�t /�  |�&/       Some_stuffs �8[�U  p9[�U  0:[justforfun_justforfun_ [�U  �<[�U  p=[�U  �=[�U  �>[�U  \�t /�  ��&/      Birthday     _Z�U  �_Z�U  �`Zjustforfun_justforfun_ Z�U  �cZ�U  `dZ�U   eZ�U  �eZ�U  ��w /�  E�&/       Meeting     �0Z�U  p1Z�U  02ZThis_stuffs_This_stuffs_ �U  �4Z�U  0?Z�U  7Z�U  �7Z�U  �/�  G5�&/      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             R�/�  r6�&/       Appointment ��[�U  @�[�U  ��[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �[�U  A�'/�  H;�&/       Birthday nt ��Z�U   �Z�U   �ZThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  `�Z�U  �̜/�  KY�&/       Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             }�/�  _�&/      Some_stuffs  �]�U  ��]�U  `�]justforfun_justforfun_ _ �U  `�]�U   �]�U  ��]�U   �]�U  �9/�  n��&/      Meeting      �Z�U  ��Z�U  `�ZThis_stuffs_This_stuffs_ �U  ��Z�U  ` [�U  `[�U   [�U  alI/�  |��&/       Workout     �^�U  `^�U  �^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �^�U   ��/�  ԧ�&/       Workout �U  ��Z�U  ��Z�U  0�ZThis_stuffs_This_stuffs_ �U  `�Z�U   �Z�U  ��Z�U  `�Z�U  ���/�  %��&/       Appointment @j]�U   k]�U  �k]justforfun_justforfun_ ]�U  �m]�U  @n]�U   o]�U  �o]�U  ���/�  s��&/      Workout     �sY�U  `tY�U  xYjustforfun_justforfun_ Y�U   �Y�U  ��Y�U  ��Y�U  ��Y�U  �a�/�  ���&/       Appointment p�Z�U  ��Z�U  ��ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p�Z�U  �q/�  )Ѩ&/      Workout     EY�U  �EY�U  �HYSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   VY�U  �/�  ���&/       Workout     �Z�U  ��Z�U   �Zjustforfun_justforfun_ Z�U  оZ�U  P�Z�U  0�Z�U  �Z�U  O�/�  !��&/      Birthday    ��X�U  ��X�U  0�XSome_stuffs_Some_stuffs_ �U   �X�U  ��X�U  ��X�U  @�X�U  �/�  `��&/       Workout                        This_stuffs_This_stuffs_                                     ��!/�  l��&/       Appointment 0�X�U  ��X�U  ��XThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��X�U  h�/�  ��&/       Appointment ��Z�U  p�Z�U  0�ZThis_stuffs_This_stuffs_ �U  ��Z�U  0�Z�U  �Z�U  ��Z�U  q��/�  ��&/       Workout     ��Y�U  @�Y�U  ��YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  � Z�U  6a�/�  �!�&/      Some_stuffs p�Y�U  0�Y�U  0�YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�Y�U  ��/�  �$�&/       Workout     0E\�U  �E\�U  PF\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  PJ\�U  ��D/�  �H�&/      Birthday    �w\�U   x\�U  �x\This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  �|\�U  $y�/�  �n�&/      Appointment 7Z�U  �7Z�U  P8Zjustforfun_justforfun_ Z�U  ;Z�U  �;Z�U  �<Z�U  P=Z�U  ��b/�  +��&/       Workout     ��Z�U  `�Z�U  ��ZThis_stuffs_This_stuffs_ �U  ��Z�U  ��Z�U  `�Z�U   �Z�U  A'n/�  ��&/       Some_stuffs 0�Z�U  �Z�U  ��ZSome_stuffs_Some_stuffs_ �U  0�Z�U  �Z�U  p�Z�U  0�Z�U  K1z/�  ��&/       Appointment 0�[�U  �[�U  p�[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��[�U  �p�/�  {��&/      Workout                        Some_stuffs_Some_stuffs_                                     -��/�  ���&/      Workout     `�^�U  ��^�U  `�^Some_stuffs_Some_stuffs_ �U  `�^�U  �^�U  `�^�U  �^�U  p /�  ���&/       Some_stuffs ��X�U  @�X�U   Yjustforfun_justforfun_ Y�U  PY�U  Y�U   	Y�U  �	Y�U  �=�/�  �&/       Workout     ��Z�U  0�Z�U  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��Z�U  �Z�/�  ��&/       Meeting �U  �Z�U  ��Z�U  p�Zjustforfun_justforfun_ Z�U  0�Z�U  ��Z�U  @�Z�U   �Z�U  
�/�  5�&/       Meeting �U  �]�U  0]�U  �]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0]�U  { �/�  {�&/       Meeting     ��\�U  p�\�U  0�\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p�\�U  �C�/�  �/�&/      Some_stuffs �cZ�U  `dZ�U   eZSome_stuffs_Some_stuffs_ �U  �gZ�U  phZ�U  0iZ�U  �iZ�U  1��/�  �1�&/       Workout ent DZ�U  �DZ�U  �EZThis_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  �IZ�U  `zp	/�  <Z�&/       Appointment ;Z�U  �;Z�U  �<ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �AZ�U  5nv	/�  �[�&/      Some_stuffs @SZ�U   TZ�U  �TZSome_stuffs_Some_stuffs_ �U  �WZ�U  @XZ�U   YZ�U  �YZ�U  �a�	/�  B|�&/       Meeting     p�\�U  0�\�U  ��\Some_stuffs_Some_stuffs_ �U  �\�U  ��\�U  p�\�U  �\�U  @O�	/�  ~�&/       Workout                        justforfun_justforfun_                                       =�	/�  7~�&/      Meeting                        justforfun_justforfun_                                       
/�  8��&/       Some_stuffs �[�U  [�U  �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  #[�U  ��
/�  L��&/       Appointment �TZ�U  �UZ�U  @VZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @[Z�U  �9�
/�  �&/      Appointment 5Y�U  �5Y�U  P8YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �EY�U  ���
/�  ���&/       Birthday    �BZ�U  PCZ�U  DZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �RZ�U  `ܭ
/�  |��&/       Appointment p�Y�U  0�Y�U  0�Yjustforfun_justforfun_ _ �U   �Y�U  ��Y�U  ��Y�U  p�Y�U  �,/�  �˪&/       Meeting ffs ��\�U   �\�U  ��\Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  �\�U  �;/�  �Ϫ&/      Appointment �[�U  ��[�U  0�[This_stuffs_This_stuffs_ �U  �[�U  p�[�U  0�[�U  ��[�U  y�D/�  Ҫ&/       Some_stuffs �\�U  ��\�U  �\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��\�U  $Z�/�  ���&/      Meeting     0�[�U  ��[�U  ��[This_stuffs_This_stuffs_ �U  ��[�U  p�[�U  0�[�U  ��[�U  x�n/�  [�&/       Appointment �l[�U   m[�U  �m[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  Pr[�U  �+q/�  �&/      Workout      D\�U  �D\�U  0E\justforfun_justforfun_ _ �U  �G\�U  PH\�U  �H\�U  PI\�U  ��x/�  � �&/       Some_stuffs  [�U  � [�U  P![This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0&[�U  0{�/�  �?�&/       Meeting     �%Y�U  �&Y�U  )YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �5Y�U  y,/�  �G�&/       Meeting     �Z�U  ��Z�U  p�Zjustforfun_justforfun_ Z�U  0�Z�U  ��Z�U  @�Z�U   �Z�U  ���/�  6i�&/       Appointment �Y�U  ��Y�U  0�YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��Y�U  ��/�  �i�&/       Meeting     p�\�U  0�\�U  ��\This_stuffs_This_stuffs_ �U  p�\�U  ��\�U  p�\�U  ��\�U  ��/�  nj�&/      Some_stuffs  �Y�U  �Y�U  0�YSome_stuffs_Some_stuffs_ �U  ��Y�U  ��Y�U  P�Y�U  �Y�U  !/�  ���&/       Birthday    p�]�U  �]�U  p�]This_stuffs_This_stuffs_ �U  p�]�U  �]�U  ��]�U  0�]�U  \�#/�  K��&/      Birthday U   �Y�U  ��Y�U  ��YSome_stuffs_Some_stuffs_ �U  P�Y�U  �Y�U  ��Y�U  ��Y�U  ˠ-/�  ͐�&/       Meeting     �y^�U  `z^�U  �z^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �~^�U  ��0/�  ���&/       Birthday     bZ�U  �bZ�U  �cZjustforfun_justforfun_ _This_stuffs_This_stuffs_ �U  phZ�U  �$�/�  ̵�&/       Birthday    ��Y�U  ��Y�U  p�YThis_stuffs_This_stuffs_ �U  ��Y�U  @�Y�U  ��Y�U  ��Y�U  ��/�  ���&/       Appointment �_]�U  ``]�U  a]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0e]�U  ��/�  P��&/      Workout     �g]�U  �h]�U  @i]Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  @m]�U  ��/�  ּ�&/       Workout     �4Z�U  0?Z�U  7ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �;Z�U  �r�/�  ���&/       Birthday     �Z�U  ��Z�U  `�ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Z�U  ��h/�  ��&/       Meeting     �Z�U  PZ�U  ZThis_stuffs_This_stuffs_ �U  `Z�U   Z�U  �Z�U  �Z�U  \�s/�  K�&/      Some_stuffs                    justforfun_justforfun_                                       u/�  ��&/       Meeting �U  0�X�U  ��X�U  ��XSome_stuffs_Some_stuffs_ �U  ��X�U  ��X�U  ��X�U  ��X�U  �M�/�  n�&/       Birthday    0_[�U  �_[�U  p`[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �d[�U  l��/�  ��&/      Appointment ��X�U  @�X�U   YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �	Y�U  Ae�/�  ��&/       Birthday    �Z�U  �%Z�U  �Zjustforfun_justforfun_ Z�U  �!Z�U  @"Z�U   #Z�U  �#Z�U  �/�  �	�&/       Meeting     puZ�U  0vZ�U  �vZThis_stuffs_This_stuffs_ �U  �yZ�U  0zZ�U  �zZ�U  �{Z�U  xf�/�  ;0�&/       Birthday     _Z�U  �_Z�U  �`ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �eZ�U  a"%/�  <S�&/       Workout      	Y�U  �	Y�U  �YThis_stuffs_This_stuffs_ �U  �Y�U  `Y�U  �Y�U  `Y�U  ��1/�  oV�&/      Appointment �Z�U  PZ�U  ZSome_stuffs_Some_stuffs_ �U  `Z�U   Z�U  �Z�U  �Z�U  �Ƽ/�  z�&/       Workout ffs  �\�U  ��\�U  @�\Some_stuffs_Some_stuffs_ �U  @�\�U   �\�U  ��\�U  ��\�U  4	�/�  �z�&/      Workout     ��X�U  @�X�U   YThis_stuffs_This_stuffs_ �U  PY�U  Y�U   	Y�U  �	Y�U  