ܦ
 /   ��
 /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �< /   �< /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     8{ /   H{ /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             | /   � /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �lw /   -mw /       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ,q /   ]q /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             \�; /   w�; /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               }f /   >}f /      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �c: /   �c: /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �|� /   /}� /   	   Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             P� /   h� /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �G- /   �G- /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             � /   9� /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��H /   ��H /      Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               l+� /   �+� /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �p� /   #q� /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �= /   �= /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                              9 /   K9 /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             4�V /   G�V /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �Ǵ /   �Ǵ /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     4� /   g� /       Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               D�v /   o�v /       Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �y /   (�y /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               X' /   p' /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               ;< /   A;< /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               � /   '� /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             -q /   ^v /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �|� /   �z� /       Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �z� /   �z� /       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ؓ� /   ٓ� /       Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             lqZ /   uqZ /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     t� /   u� /   	   Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ��� /   ��� /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             <�f /   \�f /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               �X /   �X /   	   Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     P� /   }� /       Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               N� /   $N� /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               �[, /   �[, /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��J /   ��J /   	   Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ��
 /   ��
 /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �r+ /   s+ /      Workout &V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �;i /   �;i /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��� /   N�� /       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �Г /   �Г /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     \D� /   fD� /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                                �+ /   "�+ /      Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �Ǵ /   CŴ /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             @T� /   GT� /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �*� /   �*� /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     _I /   J_I /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �TK /   �TK /       Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             du; /   �u; /      Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               h� /   �� /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     `H+ /   wH+ /   	   Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               4� /   5� /   	   Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��Z /   ��Z /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     8�w /   X�w /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �(� /   �(� /       Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               xlg /   �lg /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �|� /   Pz� /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �lw /   �ow /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             8؆ /   V؆ /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               �1 /   2 /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     4�� /   5�� /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             !9 /   9 /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             4� /   :� /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �x /   �x /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ��� /   ��� /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �lw /   �nw /   	   Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               �X /   �X /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             H�� /   {�� /   	   Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             |?� /   ~?� /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               `MX /   `MX /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     u� /   Iu� /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �: /   �: /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               m+� /   �(� /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �Y /   �Y /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             <~
 /   d~
 /      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �� /   �� /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               5� /   $� /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               <@W /   N@W /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �x /   Bx /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ��� /   ��� /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �, /   9�, /       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �-� /   �-� /      Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �1 /   . /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     � /   � /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �c: /   �f: /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ��* /   ��* /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             d� /   Fd� /      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     xO /   �O /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �r- /   �r- /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               �m� /   �m� /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             \�+ /   ��+ /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��g /   ɳg /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �p� /   dx� /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               �{h /   %|h /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �G /   D�G /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �$+ /   %+ /   	   Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��, /   ��, /       Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                              �; /   $�; /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                      �K /   <�K /       Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �+ /   "�+ /   	   Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     d� /   �� /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               0x� /   Kx� /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     u� /   6� /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               � /   �� /   	   Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �˕ /   *̕ /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��� /   ʷ� /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ��g /   ��g /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               Ԕ� /   Ք� /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     D�Z /   _�Z /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     TPu /   �Pu /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �(� /   '� /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ࡗ /   �� /       Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �h /   �h /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �
f /   �
f /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             P�K /   _�K /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ylg /   Hhg /       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �$+ /   a#+ /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �m� /   �i� /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               �[ /   �[ /   	   Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �{h /   Mwh /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �?8 /   �?8 /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ̌W /   όW /       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �� /   �� /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ��f /   ��f /       Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             8}x /   :}x /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �� /   P�� /   	   Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ��Y /   ��Y /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               ��Y /   `�Y /      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     @�w /   C�w /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               ��� /   K� /      Some_stuffs  �ҿ&V  p�ҿ&V  0��justforfun_justforfun_ ҿ&V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  ha� /   ha� /      Meeting &V  PIӿ&V  �Jӿ&V  �M�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  � /   6� /      Workout &V  ��ӿ&V  P�ӿ&V  ���justforfun_justforfun_ ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  ]�+ /   v�+ /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �p� /   �r� /      Meeting &V   �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  1x� /   �|� /      Some_stuffs PIӿ&V  �Jӿ&V  �M�justforfun_justforfun_ ӿ&V  �Vӿ&V  @Xӿ&V  p[ӿ&V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �&X /   �&X /      Birthday V  �ӿ&V  p�ӿ&V  p��Some_stuffs_Some_stuffs_ &V  �ӿ&V  `�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  L /   n /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             � X /   � X /      Appointment  �ҿ&V  p�ҿ&V  0��justforfun_justforfun_ ҿ&V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  ,�f /   >�f /      Workout &V  p[ӿ&V  �\ӿ&V  0`�justforfun_justforfun_ ӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  ��� /   ��� /   	   Appointment ��ӿ&V  p�ӿ&V  0��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  \�; /   ��; /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             !�K /   �K /       Some_stuffs  �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �� /   � /   	   Appointment PIӿ&V  �Jӿ&V  �M�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  p' /   �' /      Meeting &V  ��ӿ&V  P�ӿ&V  ���This_stuffs_This_stuffs_ &V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  D�) /   J�) /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               �uj /   �uj /       Workout &V   �ҿ&V  p�ҿ&V  0��justforfun_justforfun_ ҿ&V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  ��u /   ��u /      Some_stuffs p[ӿ&V  �\ӿ&V  0`�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  D9� /   x9� /       Birthday V  ��ӿ&V  p�ӿ&V  0��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  �5v /   �5v /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     n+� /   �"� /       Meeting &V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  ��w /   ��w /      Appointment PIӿ&V  �Jӿ&V  �M�This_stuffs_This_stuffs_ &V  �Vӿ&V  @Xӿ&V  p[ӿ&V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  � /   $� /      Some_stuffs ��ӿ&V  P�ӿ&V  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  � /   � /       Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               h�� /   ��� /      Workout &V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  ��W /   ɯW /       Workout &V  p[ӿ&V  �\ӿ&V  0`�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V   iJ /   LiJ /      Birthday V  ��ӿ&V  p�ӿ&V  0��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  �h /   ��h /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �� /   � /      Meeting &V   �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �� /   �� /       Workout &V  p[ӿ&V  �\ӿ&V  0`�justforfun_justforfun_ ӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  �� /   �� /      Some_stuffs ��ӿ&V  p�ӿ&V  0��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  �Hw /   �Hw /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �r- /   �r- /      Some_stuffs  �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �� /   W� /      Workout &V  PIӿ&V  �Jӿ&V  �M�Some_stuffs_Some_stuffs_ &V  �Vӿ&V  @Xӿ&V  p[ӿ&V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �~ /   �~ /      Appointment �ӿ&V  p�ӿ&V  p��Some_stuffs_Some_stuffs_ &V  �ӿ&V  `�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  &Z /   >&Z /      Workout &V  �6Կ&V  `8Կ&V   >�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   BԿ&V  @CԿ&V  �JԿ&V  `FԿ&V  �GԿ&V  `IԿ&V  �PԿ&V   LԿ&V  @MԿ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @      �X /   J�X /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �Z� /   �Z� /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     I�� /   ݵ� /       Appointment  �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  yO /   �S /       Appointment PIӿ&V  �Jӿ&V  �M�Some_stuffs_Some_stuffs_ &V  �Vӿ&V  @Xӿ&V  p[ӿ&V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  $>� /   8>� /      Some_stuffs �ӿ&V  p�ӿ&V  p��This_stuffs_This_stuffs_ &V  �ӿ&V  `�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  �0h /   1h /      Workout &V  �9Կ&V   ;Կ&V  �<�This_stuffs_This_stuffs_ &V  @CԿ&V  �JԿ&V  `FԿ&V  �GԿ&V  `IԿ&V  �PԿ&V   LԿ&V  @MԿ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  _I /   YI /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �� /   �� /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �� /   R� /      Meeting &V   �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  \�� /   ~�� /      Appointment PIӿ&V  �Jӿ&V  �M�Some_stuffs_Some_stuffs_ &V  �Vӿ&V  @Xӿ&V  p[ӿ&V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  Pٳ /   lٳ /      Some_stuffs ��ӿ&V  P�ӿ&V  ���This_stuffs_This_stuffs_ &V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  	&Z /   �'Z /      Appointment `FԿ&V  �GԿ&V  `I�This_stuffs_This_stuffs_ &V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  @      ��: /   ܏: /   	   Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             E�v /   ��v /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             o+� /   �(� /      Some_stuffs  �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �ky /   �ky /       Meeting     �Vӿ&V  @Xӿ&V  p[�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  �� /   �� /      Meeting &V  ��ӿ&V  P�ӿ&V  ���Some_stuffs_Some_stuffs_ &V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  AT� /   W� /       Workout &V  `IԿ&V  �PԿ&V   L�justforfun_justforfun_ Կ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  pԿ&V  �xԿ&V  �� /   ¤ /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     i� /   � /      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     <GZ /   cGZ /      Appointment  �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �[ /   �[ /      Some_stuffs p[ӿ&V  �\ӿ&V  0`�justforfun_justforfun_ ӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  L�h /   �h /       Some_stuffs ��ӿ&V  p�ӿ&V  0��This_stuffs_This_stuffs_ &V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  @b� /   ub� /      Meeting &V   RԿ&V  �SԿ&V   U�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  pԿ&V  �xԿ&V  �yԿ&V  p{Կ&V  �|Կ&V  ��Կ&V   �Կ&V  ��Կ&V  �^� /   �^� /      Meeting &V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V   /   E /      Appointment p[ӿ&V  �\ӿ&V  0`�This_stuffs_This_stuffs_ &V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  �H /    �H /      Appointment ��ӿ&V  p�ӿ&V  0��This_stuffs_This_stuffs_ &V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  �G /   x�G /      Appointment  RԿ&V  �SԿ&V   U�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  pԿ&V  �xԿ&V  �yԿ&V  p{Կ&V  �|Կ&V  ��Կ&V   �Կ&V  ��Կ&V  |�* /   ��* /      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ��8 /   ��8 /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               � /   � /   	   Appointment  �ҿ&V  p�ҿ&V  0��justforfun_justforfun_ ҿ&V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  ]�� /   4�� /      Some_stuffs PIӿ&V  �Jӿ&V  �M�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �؈ /   �؈ /   	   Meeting &V  �ӿ&V  p�ӿ&V  p��This_stuffs_This_stuffs_ &V  �ӿ&V  `�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  � /   �� /      Birthday V  �9Կ&V   ;Կ&V  �<�justforfun_justforfun_ Կ&V  @CԿ&V  �JԿ&V  `FԿ&V  �GԿ&V  `IԿ&V  �PԿ&V   LԿ&V  @MԿ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  �� /   �� /   	   Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     <1f /   Q1f /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     u� /   Qo� /      Workout &V   �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  M�h /   ��h /      Meeting     PIӿ&V  �Jӿ&V  �M�Some_stuffs_Some_stuffs_ &V  �Vӿ&V  @Xӿ&V  p[ӿ&V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �� /   � /      Birthday V  �ӿ&V  p�ӿ&V  p��justforfun_justforfun_ ӿ&V  �ӿ&V  `�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  �� /   � /      Birthday V  �9Կ&V   ;Կ&V  �<�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �GԿ&V  `IԿ&V  �PԿ&V   LԿ&V  @MԿ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  �[, /   (^, /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             A�w /   ��w /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �Г /   �ԓ /   	   Appointment  �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  ��H /   ��H /      Workout     PIӿ&V  �Jӿ&V  �M�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �
f /   �f /   	   Meeting     �ӿ&V  p�ӿ&V  p��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  P�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  0) /   _) /      Meeting &V  �(Կ&V  P*Կ&V  �/�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   ;Կ&V  �<Կ&V   EԿ&V  �@Կ&V   BԿ&V  @CԿ&V  �JԿ&V  `FԿ&V  �GԿ&V  `IԿ&V  �PԿ&V   LԿ&V  @MԿ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  �̲ /   Ͳ /      Workout &V  `sԿ&V  �tԿ&V  0~�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   �Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  @�Կ&V  @�Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  `�Կ&V  0�Կ&V  p�Կ&V   �Կ&V  @�Կ&V  ��Կ&V   �Կ&V  P�Կ&V  ��Կ&V  �Կ&V  0�Կ&V  p�Կ&V  ,�< /   P�< /      Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �� /   �� /      Birthday V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  ��f /   ȣf /      Appointment p[ӿ&V  �\ӿ&V  0`�justforfun_justforfun_ ӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  �5* /   �5* /      Some_stuffs ��ӿ&V  P�ӿ&V  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  H�� /   K�� /      Birthday V  `FԿ&V  �GԿ&V  `I�Some_stuffs_Some_stuffs_ &V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  ��9 /   ��9 /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     }�* /   q�* /       Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               PPj /   gPj /      Birthday V   �ҿ&V  p�ҿ&V  0��justforfun_justforfun_ ҿ&V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �� /   /� /   	   Some_stuffs p[ӿ&V  �\ӿ&V  0`�Some_stuffs_Some_stuffs_ &V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  X=� /   p=� /      Birthday    ��ӿ&V  P�ӿ&V  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  �� /   �� /      Workout &V  `FԿ&V  �GԿ&V  `I�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  ᡗ /   E�� /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               � X /   ��W /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     E�Z /   ��Z /       Birthday V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  � /   ȥ /       Birthday    PIӿ&V  �Jӿ&V  �M�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �� /   m�� /   	   Birthday    �ӿ&V  `�ӿ&V  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V   �� /   �� /      Birthday V   >Կ&V  @?Կ&V  �9�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �JԿ&V  `FԿ&V  �GԿ&V  `IԿ&V  �PԿ&V   LԿ&V  @MԿ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  Y=� /   :;� /      Birthday V  0~Կ&V  pԿ&V  �x�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  `�Կ&V  ��Կ&V  @�Կ&V  @�Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  `�Կ&V  0�Կ&V  p�Կ&V   �Կ&V  @�Կ&V  ��Կ&V   �Կ&V  P�Կ&V  ��Կ&V  �Կ&V  0�Կ&V  p�Կ&V  �Կ&V  `�Կ&V  �x /   �x /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �m� /   �m� /      Workout &V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  ��g /   ��g /      Meeting     p[ӿ&V  �\ӿ&V  0`�This_stuffs_This_stuffs_ &V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  X�� /   f�� /      Appointment ��ӿ&V  p�ӿ&V  0��This_stuffs_This_stuffs_ &V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  �� /   @� /      Birthday V   RԿ&V  �SԿ&V   U�justforfun_justforfun_ Կ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  pԿ&V  �xԿ&V  �yԿ&V  p{Կ&V  �|Կ&V  ��Կ&V   �Կ&V  ��Կ&V  l$� /   �$� /      Meeting &V  `�Կ&V  ��Կ&V  `��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  p�Կ&V   �Կ&V  @�Կ&V  ��Կ&V   �Կ&V  P�Կ&V  ��Կ&V  �Կ&V  0�Կ&V  p�Կ&V  �Կ&V  `�Կ&V  ��Կ&V  ЩԿ&V  �Կ&V  P�Կ&V  ��Կ&V  �Կ&V  ��Կ&V  �Կ&V  `�Կ&V  ��Կ&V   �Կ&V  ��Կ&V  �Կ&V  �Կ&V  �r- /   Wq- /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             в� /   㲖 /      Meeting &V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �_� /   �_� /       Appointment p[ӿ&V  �\ӿ&V  0`�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  e� /   K� /      Appointment ��ӿ&V  p�ӿ&V  0��This_stuffs_This_stuffs_ &V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  !�; /   q�; /      Some_stuffs `FԿ&V  �GԿ&V  `I�justforfun_justforfun_ Կ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  8�I /   :�I /      Appointment ��Կ&V   �Կ&V  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  ��Կ&V  `�Կ&V  ��Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  `�Կ&V  0�Կ&V  p�Կ&V   �Կ&V  @�Կ&V  ��Կ&V   �Կ&V  P�Կ&V  ��Կ&V  �Կ&V  0�Կ&V  p�Կ&V  �Կ&V  `�Կ&V  ��Կ&V  ЩԿ&V  �Կ&V  P�Կ&V  ��Կ&V  �Կ&V  �H /   ��H /   	   Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �^< /   �^< /      Birthday V   �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  0O� /   :O� /      Appointment p[ӿ&V  �\ӿ&V  0`�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  hH /   �H /      Appointment ��ӿ&V  p�ӿ&V  0��This_stuffs_This_stuffs_ &V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  Dף /   wף /      Workout &V   RԿ&V  �SԿ&V   U�Some_stuffs_Some_stuffs_ &V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  pԿ&V  �xԿ&V  �yԿ&V  p{Կ&V  �|Կ&V  ��Կ&V   �Կ&V  ��Կ&V  ݦ
 /   ��
 /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �< /   �< /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     9{ /   H{ /      Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  } /   � /      Workout     P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �lw /   -mw /       Some_stuffs ��/V  p�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  .q /   ]q /      Some_stuffs  ��/V  @��/V  ��Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ]�; /   w�; /      Meeting /V  ���/V   ��/V  `�justforfun_justforfun_ �/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  }f /   >}f /      Workout /V  �	�/V  �/V  PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �c: /   �c: /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �|� /   /}� /   	   Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             Q� /   h� /      Birthday V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �G- /   �G- /      Meeting     P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  � /   9� /      Some_stuffs ��/V  p�/V  pThis_stuffs_This_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  ��H /   ��H /      Some_stuffs Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  p+� /   �+� /      Some_stuffs ���/V  ���/V   �Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  �p� /   #q� /      Birthday V  � �/V  0�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  �= /   �= /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             "9 /   K9 /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             5�V /   G�V /      Birthday V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �Ǵ /   �Ǵ /      Birthday    P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  5� /   g� /       Birthday    ��/V  p�/V  pjustforfun_justforfun_ �/V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  F�v /   o�v /       Workout     Ј�/V  P��/V  ЏThis_stuffs_This_stuffs_ /V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  �y /   (�y /      Workout /V  ���/V  ���/V   �justforfun_justforfun_ �/V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  Y' /   p' /      Birthday V  � �/V  0�/V  pjustforfun_justforfun_ �/V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  ;< /   A;< /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               � /   '� /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             /q /   ^v /      Birthday V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �|� /   �z� /       Some_stuffs ���/V  @��/V  p�Some_stuffs_Some_stuffs_ /V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  �z� /   �z� /       Workout     ��/V  `�/V  �#Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  ٓ� /   ٓ� /       Some_stuffs  ��/V  @��/V  ��This_stuffs_This_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  mqZ /   uqZ /      Meeting /V  ���/V   ��/V  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  v� /   u� /   	   Workout /V  �	�/V  �/V  PSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  ��� /   ��� /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             =�f /   \�f /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               �X /   �X /   	   Some_stuffs  U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  Q� /   }� /       Some_stuffs P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  N� /   $N� /      Appointment ��/V  p�/V  pjustforfun_justforfun_ �/V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  �[, /   �[, /      Birthday    Ј�/V  P��/V  ЏThis_stuffs_This_stuffs_ /V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  ��J /   ��J /   	   Meeting /V  ���/V  ���/V   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  ��
 /   ��
 /      Some_stuffs � �/V  0�/V  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  �r+ /   s+ /      Workout /V   <�/V  �F�/V  @?This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  �;i /   �;i /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��� /   N�� /       Some_stuffs  U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �Г /   �Г /      Workout     ���/V  @��/V  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  ]D� /   fD� /      Meeting     ��/V  `�/V  �#justforfun_justforfun_ �/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  �+ /   "�+ /      Appointment  ��/V  @��/V  ��This_stuffs_This_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  �Ǵ /   CŴ /      Some_stuffs ���/V   ��/V  `�Some_stuffs_Some_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  BT� /   GT� /      Birthday V  ��/V  `�/V  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  �*� /   �*� /      Birthday V  `M�/V  �N�/V  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  @      _I /   J_I /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �TK /   �TK /       Appointment  U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  eu; /   �u; /      Some_stuffs P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  j� /   �� /      Workout     ��/V  p�/V  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  aH+ /   wH+ /   	   Some_stuffs Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  6� /   5� /   	   Some_stuffs ���/V  ���/V   �This_stuffs_This_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  ��Z /   ��Z /      Some_stuffs � �/V  0�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  9�w /   X�w /      Some_stuffs  <�/V  �F�/V  @?Some_stuffs_Some_stuffs_ /V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  �(� /   �(� /       Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               zlg /   �lg /      Workout /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �|� /   Pz� /      Workout     P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �lw /   �ow /      Some_stuffs ��/V  p�/V  pSome_stuffs_Some_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  9؆ /   V؆ /      Appointment Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  �1 /   2 /      Appointment ���/V  ���/V   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  5�� /   5�� /      Meeting /V  � �/V  0�/V  pThis_stuffs_This_stuffs_ /V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  #9 /   9 /      Birthday V   <�/V  �F�/V  @?Some_stuffs_Some_stuffs_ /V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  5� /   :� /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �x /   �x /      Workout /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ��� /   ��� /      Some_stuffs P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �lw /   �nw /   	   Some_stuffs ��/V  p�/V  pjustforfun_justforfun_ �/V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  �X /   �X /      Some_stuffs ���/V   ��/V  ��Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  J�� /   {�� /   	   Workout     p��/V  ���/V  ��Some_stuffs_Some_stuffs_ /V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �/V  P�/V  }?� /   ~?� /      Meeting /V  ��/V   �/V  �!justforfun_justforfun_ �/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  aMX /   `MX /      Meeting /V  �Z�/V  �[�/V  �RSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V  u� /   Iu� /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �: /   �: /      Birthday V   U�/V  pW�/V  0Yjustforfun_justforfun_ �/V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  q+� /   �(� /      Meeting     P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �Y /   �Y /      Workout     �#�/V  P%�/V  �)This_stuffs_This_stuffs_ /V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  =~
 /   d~
 /      Workout     ���/V   ��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  �� /   �� /      Workout     `��/V  ���/V  0�justforfun_justforfun_ �/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  7� /   $� /      Birthday V  P�/V  ��/V  justforfun_justforfun_ �/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  =@W /   N@W /      Appointment �Z�/V  �[�/V  �RSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V  �x /   Bx /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ��� /   ��� /      Some_stuffs  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �, /   9�, /       Meeting     P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �-� /   �-� /      Appointment ��/V  p�/V  pThis_stuffs_This_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  �1 /   . /      Workout     Ј�/V  P��/V  ЏSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  � /   � /      Birthday    ���/V   ��/V  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  �c: /   �f: /      Appointment �	�/V  �/V  PSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  ��* /   ��* /      Some_stuffs `M�/V  �N�/V  �ZSome_stuffs_Some_stuffs_ /V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  d� /   Fd� /      Workout /V  ���/V  0��/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  @      zO /   �O /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �r- /   �r- /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               �m� /   �m� /      Some_stuffs  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ^�+ /   ��+ /      Birthday    P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��g /   ɳg /      Workout     ��/V  p�/V  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  �p� /   dx� /      Appointment Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  �{h /   %|h /      Workout     ���/V  ���/V   �Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  �G /   D�G /      Appointment � �/V  0�/V  pSome_stuffs_Some_stuffs_ /V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  �$+ /   %+ /   	   Meeting /V   <�/V  �F�/V  @?Some_stuffs_Some_stuffs_ /V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  ��, /   ��, /       Meeting /V  0s�/V  pt�/V  �uThis_stuffs_This_stuffs_ /V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  "�; /   $�; /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     "�K /   <�K /       Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �+ /   "�+ /   	   Meeting /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  f� /   �� /      Birthday    ���/V  @��/V  p�justforfun_justforfun_ �/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  2x� /   Kx� /      Birthday    ��/V  `�/V  �#This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  w� /   6� /      Birthday     ��/V  @��/V  ��justforfun_justforfun_ �/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  � /   �� /   	   Workout     ���/V  ���/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �˕ /   *̕ /      Meeting     ��/V   �/V  p+This_stuffs_This_stuffs_ /V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  ��� /   ʷ� /      Meeting /V  �W�/V  �X�/V  �eSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  ��g /   ��g /      Appointment ���/V  0��/V  p�justforfun_justforfun_ �/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  Ք� /   Ք� /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     F�Z /   _�Z /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     UPu /   �Pu /      Appointment  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �(� /   '� /      Birthday    P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ⡗ /   �� /       Appointment ��/V  p�/V  pSome_stuffs_Some_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  �h /   �h /      Birthday    Ј�/V  P��/V  ЏSome_stuffs_Some_stuffs_ /V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  �
f /   �
f /      Birthday    ���/V  ���/V   �Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  Q�K /   _�K /      Some_stuffs � �/V  0�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  {lg /   Hhg /       Meeting /V   <�/V  �F�/V  @?Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  �$+ /   a#+ /      Meeting /V  �z�/V  ���/V  �~Some_stuffs_Some_stuffs_ /V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  �m� /   �i� /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               �[ /   �[ /   	   Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �{h /   Mwh /      Meeting /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �?8 /   �?8 /      Some_stuffs ���/V  @��/V  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  ͌W /   όW /       Meeting     ��/V  `�/V  �#Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  �� /   �� /      Meeting      ��/V  @��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ��f /   ��f /       Appointment ���/V   ��/V  `�Some_stuffs_Some_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  9}x /   :}x /      Meeting     �	�/V  �/V  PThis_stuffs_This_stuffs_ /V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �� /   P�� /   	   Appointment P�/V  PQ�/V  0HThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  ��Y /   ��Y /      Appointment �z�/V  ���/V  �~justforfun_justforfun_ �/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  ��Y /   `�Y /      Appointment ���/V  P��/V  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V  B�w /   C�w /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               ��� /   K� /      Some_stuffs  U�/V  pW�/V  0Yjustforfun_justforfun_ �/V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ia� /   ha� /      Meeting     ���/V  @��/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  � /   6� /      Workout     ��/V  `�/V  �#justforfun_justforfun_ �/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  _�+ /   v�+ /      Workout      ��/V  @��/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  �p� /   �r� /      Meeting     ���/V  ���/V  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  3x� /   �|� /      Some_stuffs ��/V  `�/V  �justforfun_justforfun_ �/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  �&X /   �&X /      Birthday V  U�/V  PV�/V  �WSome_stuffs_Some_stuffs_ /V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  M /   n /      Meeting /V  p��/V  ���/V  ��This_stuffs_This_stuffs_ /V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  � X /   � X /      Appointment ���/V  ���/V  �justforfun_justforfun_ �/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  -�f /   >�f /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               ��� /   ��� /   	   Appointment  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ]�; /   ��; /      Workout     P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  #�K /   �K /       Some_stuffs ��/V  p�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  �� /   � /   	   Appointment  ��/V  @��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  q' /   �' /      Meeting     ���/V   ��/V  `�This_stuffs_This_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  E�) /   J�) /      Meeting     �	�/V  �/V  Pjustforfun_justforfun_ �/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �uj /   �uj /       Workout     P�/V  PQ�/V  0Hjustforfun_justforfun_ �/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  ��u /   ��u /      Some_stuffs �z�/V  ���/V  �~This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  E9� /   x9� /       Birthday V  ���/V  P��/V  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V  �5v /   �5v /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     r+� /   �"� /       Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ��w /   ��w /      Appointment P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  � /   $� /      Some_stuffs ��/V  p�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  � /   � /       Some_stuffs Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  i�� /   ��� /      Workout     ���/V   ��/V  `�This_stuffs_This_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  ��W /   ɯW /       Workout     �	�/V  �/V  PSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  !iJ /   LiJ /      Birthday    P�/V  PQ�/V  0HThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  �h /   ��h /      Meeting /V  �z�/V  ���/V  �~This_stuffs_This_stuffs_ /V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  �� /   � /      Meeting /V   ��/V  `��/V  мSome_stuffs_Some_stuffs_ /V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  �� /   �� /       Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               �� /   �� /      Some_stuffs  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �Hw /   �Hw /      Meeting     ���/V  @��/V  p�Some_stuffs_Some_stuffs_ /V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  �r- /   �r- /      Some_stuffs ��/V  `�/V  �#Some_stuffs_Some_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  �� /   W� /      Workout      ��/V  @��/V  ��Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  �~ /   �~ /      Appointment ���/V   ��/V  `�Some_stuffs_Some_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  
&Z /   >&Z /      Workout     �	�/V  �/V  PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �X /   J�X /      Workout     P�/V  PQ�/V  0HSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  �Z� /   �Z� /      Appointment �z�/V  ���/V  �~Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  K�� /   ݵ� /       Appointment ���/V  P��/V  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V  {O /   �S /       Appointment @��/V  ���/V  ��Some_stuffs_Some_stuffs_ /V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @      %>� /   8>� /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �0h /   1h /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             _I /   YI /      Birthday V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �� /   �� /      Workout     ���/V  @��/V  p�Some_stuffs_Some_stuffs_ /V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  �� /   R� /      Meeting     ��/V  `�/V  �#Some_stuffs_Some_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  ^�� /   ~�� /      Appointment @��/V  ���/V  `�Some_stuffs_Some_stuffs_ /V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  `��/V  0��/V  p��/V  ���/V   ��/V  `��/V  Qٳ /   lٳ /      Some_stuffs p��/V  ���/V  ��This_stuffs_This_stuffs_ /V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �/V  P�/V  &Z /   �'Z /      Appointment ��/V   �/V  �!This_stuffs_This_stuffs_ /V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  ��: /   ܏: /   	   Some_stuffs �W�/V  �X�/V  �eThis_stuffs_This_stuffs_ /V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  G�v /   ��v /      Appointment ���/V  0��/V  p�Some_stuffs_Some_stuffs_ /V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  s+� /   �(� /      Some_stuffs ���/V   ��/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V  �ky /   �ky /       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �� /   �� /      Meeting /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  CT� /   W� /       Workout     P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �� /   ¤ /      Some_stuffs ��/V  `�/V  �#Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  k� /   � /      Workout      ��/V  @��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  =GZ /   cGZ /      Appointment ���/V  ���/V  p�This_stuffs_This_stuffs_ /V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �[ /   �[ /      Some_stuffs ��/V  `�/V  �justforfun_justforfun_ �/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  N�h /   �h /       Some_stuffs `M�/V  �N�/V  �ZThis_stuffs_This_stuffs_ /V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  Ab� /   ub� /      Meeting     ���/V  0��/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  �^� /   �^� /      Meeting /V   ��/V  `��/V  мThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V   /   E /      Appointment @��/V  ���/V  ��This_stuffs_This_stuffs_ /V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �H /    �H /      Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �G /   x�G /      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ~�* /   ��* /      Appointment  U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ��8 /   ��8 /      Meeting     P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  � /   � /   	   Appointment ��/V  p�/V  pjustforfun_justforfun_ �/V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  _�� /   4�� /      Some_stuffs Ј�/V  P��/V  ЏThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  �؈ /   �؈ /   	   Meeting     ���/V   ��/V  `�This_stuffs_This_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  � /   �� /      Birthday    �	�/V  �/V  Pjustforfun_justforfun_ �/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �� /   �� /   	   Workout     P�/V  PQ�/V  0HSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  =1f /   Q1f /      Some_stuffs �z�/V  ���/V  �~Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  u� /   Qo� /      Workout /V  ���/V  P��/V  �Some_stuffs_Some_stuffs_ /V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V  O�h /   ��h /      Meeting /V  @��/V  ���/V  ��Some_stuffs_Some_stuffs_ /V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �� /   � /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �� /   � /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �[, /   (^, /      Some_stuffs  U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  C�w /   ��w /      Appointment P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �Г /   �ԓ /   	   Appointment ��/V  `�/V  �#This_stuffs_This_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  ��H /   ��H /      Workout     ���/V   ��/V  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  `��/V  0��/V  p��/V  ���/V  �
f /   �f /   	   Meeting     ���/V  `��/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  1) /   _) /      Meeting     P$�/V  �%�/V   'This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  �̲ /   Ͳ /      Workout     0]�/V  p^�/V  �_This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  -�< /   P�< /      Appointment ���/V  Д�/V  �This_stuffs_This_stuffs_ /V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  �� /   �� /      Birthday V  ��/V  P��/V  ��This_stuffs_This_stuffs_ /V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ��f /   ȣf /      Appointment @��/V  � 	�/V  �	justforfun_justforfun_ 	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  �5* /   �5* /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     I�� /   K�� /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��9 /   ��9 /      Meeting /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �* /   q�* /       Meeting     P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  QPj /   gPj /      Birthday    ��/V  `�/V  �#justforfun_justforfun_ �/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  �� /   /� /   	   Some_stuffs  ��/V  @��/V  ��Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  Z=� /   p=� /      Birthday    ���/V  ���/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �� /   �� /      Workout     ��/V  `�/V  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  㡗 /   E�� /      Workout     `M�/V  �N�/V  �Zjustforfun_justforfun_ �/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  � X /   ��W /      Meeting     p��/V  ���/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  G�Z /   ��Z /       Birthday V  ��/V  P��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  � /   ȥ /       Birthday V  �	�/V  P	�/V  �		This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �� /   m�� /   	   Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �� /   �� /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     [=� /   :;� /      Birthday V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �x /   �x /      Birthday    ���/V  @��/V  p�This_stuffs_This_stuffs_ /V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  �m� /   �m� /      Workout     ��/V  `�/V  �#This_stuffs_This_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  ��g /   ��g /      Meeting      ��/V  @��/V  ��This_stuffs_This_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  Y�� /   f�� /      Appointment ���/V   ��/V  `�This_stuffs_This_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  �� /   @� /      Birthday    �	�/V  �/V  Pjustforfun_justforfun_ �/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  m$� /   �$� /      Meeting     �Z�/V  �[�/V  �RSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V  �r- /   Wq- /      Meeting     p��/V  P��/V  ��This_stuffs_This_stuffs_ /V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  Ѳ� /   㲖 /      Meeting     м�/V  ��/V  @�This_stuffs_This_stuffs_ /V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  �_� /   �_� /       Appointment ���/V   ��/V  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V  g� /   K� /      Appointment `'	�/V  �(	�/V  �)	This_stuffs_This_stuffs_ /V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  �R	�/V  T	�/V  #�; /   q�; /      Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               9�I /   :�I /      Appointment  U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �H /   ��H /   	   Meeting     P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �^< /   �^< /      Birthday    ��/V  `�/V  �#Some_stuffs_Some_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  1O� /   :O� /      Appointment  ��/V  @��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  iH /   �H /      Appointment ���/V   ��/V  `�This_stuffs_This_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  Eף /   wף /      Workout     �	�/V  �/V  PSome_stuffs_Some_stuffs_ /V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �-� /   n1� /      Meeting     P�/V  PQ�/V  0HSome_stuffs_Some_stuffs_ /V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  >~
 /   �}
 /      Appointment �z�/V  ���/V  �~This_stuffs_This_stuffs_ /V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  lŗ /   �ŗ /      Birthday    ���/V  P��/V  �This_stuffs_This_stuffs_ /V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V  �t) /   �t) /      Workout     ���/V  ���/V  �Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  P� /   �� /      Workout /V  @	�/V  �,	�/V  �	justforfun_justforfun_ 	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  h� /   �� /      Meeting /V  �Q	�/V  �R	�/V  T	Some_stuffs_Some_stuffs_ /V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  �|� /   �x� /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               L�V /   l�V /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               2) /   k) /      Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �Г /   qՓ /      Appointment P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �x /   �x /      Birthday    ��/V  p�/V  pSome_stuffs_Some_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  N /   � /       Birthday    Ј�/V  P��/V  ЏThis_stuffs_This_stuffs_ /V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  d� /   e� /      Appointment ���/V  ���/V   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  w /   "w /      Birthday    � �/V  0�/V  pjustforfun_justforfun_ �/V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  �X /   ��X /      Appointment  <�/V  �F�/V  @?Some_stuffs_Some_stuffs_ /V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   R9 /   /R9 /      Appointment 0s�/V  pt�/V  �uSome_stuffs_Some_stuffs_ /V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  |D /   �D /      Appointment ���/V  Ъ�/V  P�justforfun_justforfun_ �/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V  >@W /   -AW /      Some_stuffs ���/V   ��/V  @�Some_stuffs_Some_stuffs_ /V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  XaG /   �aG /      Birthday V  `	�/V  �	�/V  	This_stuffs_This_stuffs_ /V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  ��� /   ã� /   	   Birthday V  PZ	�/V  �[	�/V  `L	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �H /   <�H /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             :�w /   q�w /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ~ /   f /      Workout /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V    /   Y /      Workout     P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  Rٳ /   �۳ /      Birthday    ��/V  p�/V  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  p�Y /   ��Y /      Meeting     Ј�/V  P��/V  ЏSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V   /    /      Workout     ���/V  ���/V   �This_stuffs_This_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  �� /   � /      Meeting     � �/V  0�/V  pThis_stuffs_This_stuffs_ /V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  dW /   �W /      Meeting      <�/V  �F�/V  @?Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  >1f /   /f /      Meeting     0s�/V  pt�/V  �uThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  &>� /   �>� /      Meeting     ���/V  Ъ�/V  P�justforfun_justforfun_ �/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V  4�v /   X�v /      Appointment ���/V   ��/V  @�This_stuffs_This_stuffs_ /V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  h /   h /      Meeting /V  `	�/V  �	�/V  	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  Н) /   ��) /      Birthday V  PZ	�/V  �[	�/V  `L	This_stuffs_This_stuffs_ /V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  T~� /   W~� /       Appointment ��	�/V  ��	�/V   �	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  ?1f /   �1f /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     4�� /   4�� /      Some_stuffs  U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ��g /   ��g /      Some_stuffs P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  :�I /   ��I /       Some_stuffs ��/V  p�/V  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  ��i /   ��i /      Meeting     Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  	 /   _ /      Workout     ���/V  ���/V   �Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  � /   �� /      Meeting     � �/V  0�/V  pjustforfun_justforfun_ �/V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  �$+ /   �"+ /      Meeting      <�/V  �F�/V  @?justforfun_justforfun_ �/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  eW /   �W /      Meeting     0s�/V  pt�/V  �uThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  Q� /   Q� /      Birthday    ���/V  Ъ�/V  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V  ģ9 /   ��9 /      Meeting     ���/V   ��/V  @�justforfun_justforfun_ �/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  !R9 /   �W9 /      Meeting     `	�/V  �	�/V  	This_stuffs_This_stuffs_ /V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  Z' /   �* /      Birthday V  PZ	�/V  �[	�/V  `L	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �+ /   �+ /   	   Meeting /V  ��	�/V  ��	�/V   �	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  �� /   �� /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �
f /   �	f /      Some_stuffs  U�/V  pW�/V  0Yjustforfun_justforfun_ �/V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �X /   5�X /      Appointment P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �2I /   �2I /      Appointment ��/V  `�/V  �#This_stuffs_This_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  $ /   [ /      Birthday     ��/V  @��/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  �<Y /   �<Y /   	   Appointment ���/V   ��/V  `�Some_stuffs_Some_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  �� /   >�� /      Birthday    �	�/V  �/V  PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �[ /   7[ /      Appointment P�/V  PQ�/V  0HSome_stuffs_Some_stuffs_ /V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  �j� /   �j� /       Appointment �z�/V  ���/V  �~Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  $9 /   l9 /      Appointment ���/V  P��/V  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V  O /   ) /   	   Appointment ���/V  ���/V  �Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �TK /   �SK /       Workout     �$	�/V   &	�/V  `'	Some_stuffs_Some_stuffs_ /V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  ��f /   x�f /   	   Some_stuffs  k	�/V  `l	�/V  �\	Some_stuffs_Some_stuffs_ /V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V   �	�/V  @�	�/V  \U; /   �U; /      Workout /V  �	�/V  P�	�/V  ��	This_stuffs_This_stuffs_ /V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  Ю	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  fW /   �W /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             $�v /   K�v /      Workout /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �5v /   �8v /       Birthday    p��/V  ��/V  0�This_stuffs_This_stuffs_ /V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  p�/V  p�/V  >GZ /   �HZ /      Appointment �#�/V  P%�/V  �)This_stuffs_This_stuffs_ /V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  p� /   �� /      Appointment ���/V   ��/V  ��Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  �� /   �� /   	   Appointment ���/V   ��/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �/V  P�/V  ��/V  �/V  0q /   3p /      Appointment P$�/V  �%�/V   'justforfun_justforfun_ �/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  ��9 /   *�9 /      Workout     0]�/V  p^�/V  �_This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ��u /   ��u /       Some_stuffs ���/V  Д�/V  �justforfun_justforfun_ �/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  (�J /   <�J /      Appointment  ��/V  ���/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  Hu� /   ou� /      Appointment `	�/V  �	�/V  	Some_stuffs_Some_stuffs_ /V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  HBg /   {Bg /      Birthday V  T	�/V  PU	�/V  �V	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  6� /   � /      Appointment �	�/V  P�	�/V  ��	This_stuffs_This_stuffs_ /V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  Ю	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  �Y /   �Y /   	   Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �� /   7�� /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               �� /   �� /      Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ! /   A /      Appointment p��/V  ��/V  0�justforfun_justforfun_ �/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  p�/V  p�/V  �;� /   �;� /      Appointment �#�/V  P%�/V  �)Some_stuffs_Some_stuffs_ /V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  fu; /   �u; /      Appointment `��/V  ��/V  `�This_stuffs_This_stuffs_ /V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  `��/V  0��/V  p��/V  ���/V   ��/V  `��/V  ���/V  0��/V  q� /   �� /   	   Some_stuffs ���/V   ��/V  ��Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �/V  P�/V  ��/V  �/V  �Q /   R /      Workout     �!�/V  #�/V  �Some_stuffs_Some_stuffs_ /V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V  ��8 /   /�8 /      Appointment 0]�/V  p^�/V  �_justforfun_justforfun_ �/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  t�i /   ~�i /      Appointment ���/V  Д�/V  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  gi /   gi /      Appointment  ��/V  ���/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  _v /   1_v /      Appointment `	�/V  �	�/V  	Some_stuffs_Some_stuffs_ /V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  �E� /   �E� /      Some_stuffs T	�/V  PU	�/V  �V	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  0ou /   Jou /      Some_stuffs �	�/V  P�	�/V  ��	Some_stuffs_Some_stuffs_ /V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  Ю	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��x /   �x /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               �Y /    Y /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �< /   E< /       Workout /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �< /   �< /      Workout     P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �� /   �� /      Appointment ��/V  `�/V  �#This_stuffs_This_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  �: /   �: /       Birthday     ��/V  @��/V  ��This_stuffs_This_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  �y /   �y /      Some_stuffs ���/V   ��/V  `�justforfun_justforfun_ �/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  �+ /   )�+ /   	   Birthday    ��/V   �/V  �!justforfun_justforfun_ �/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  �Q /   "R /      Birthday    �e�/V  �f�/V  0]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  �Q /   4N /      Workout     p��/V  0��/V  ��Some_stuffs_Some_stuffs_ /V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ��
 /   k�
 /      Some_stuffs ���/V  ���/V  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V  �+ /   Ù+ /      Meeting     ���/V  ���/V  @�justforfun_justforfun_ 	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  �$+ /   $+ /      Workout     �0	�/V   2	�/V  @3	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  "J /   -"J /      Meeting     �g	�/V  �h	�/V  P|	This_stuffs_This_stuffs_ /V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  h�< /   ��< /      Appointment ��	�/V  Щ	�/V  �	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  C /   6C /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     }f /   {}f /      Workout /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  D�w /   8�w /      Appointment P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �� /   7� /      Workout     ��/V  p�/V  pThis_stuffs_This_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  6�V /   ��V /      Birthday    Ј�/V  P��/V  ЏThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  p�I /   ��I /      Birthday    ���/V  ���/V   �This_stuffs_This_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  ��� /   ��� /      Birthday    P�/V  ��/V  Some_stuffs_Some_stuffs_ /V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  ��Z /   ��Z /      Meeting     �R�/V  �S�/V  UThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ԨG /   �G /      Birthday    ���/V  0��/V  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ��� /   ��� /   	   Workout     ��/V  P��/V  ��This_stuffs_This_stuffs_ /V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  �� /   �� /      Birthday    �		�/V  �
	�/V  	Some_stuffs_Some_stuffs_ /V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  �� /   W� /       Birthday    PZ	�/V  �[	�/V  `L	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �P� /   �P� /      Appointment ��	�/V  ��	�/V   �	Some_stuffs_Some_stuffs_ /V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  X�� /   n�� /      Some_stuffs �	�/V  0�	�/V  p�	Some_stuffs_Some_stuffs_ /V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  p�	�/V  @�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V   �	�/V  `�	�/V  ��	�/V  P�	�/V  ��	�/V  0�	�/V  p�	�/V  � /   �� /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               r' /   K( /      Appointment  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  h-9 /   p-9 /   	   Birthday    P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �A� /   B� /      Workout     �#�/V  P%�/V  �)Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  ��( /   ��( /      Meeting     `��/V  ��/V  `�justforfun_justforfun_ �/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  `��/V  0��/V  p��/V  ���/V   ��/V  `��/V  ���/V  0��/V  䡗 /   )�� /   	   Some_stuffs `��/V  ���/V  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  ��W /   d�W /      Appointment P$�/V  �%�/V   'This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  u� /   =o� /      Appointment 0]�/V  p^�/V  �_Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ^�; /   ��; /      Appointment ���/V  Д�/V  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ��X /   \�X /      Some_stuffs ��/V  P��/V  ��justforfun_justforfun_ �/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  �˕ /   
ʕ /      Appointment @��/V  � 	�/V  �	This_stuffs_This_stuffs_ /V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  �+ /   �+ /      Workout     @3	�/V  �4	�/V  �5	justforfun_justforfun_ 	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �{h /   &xh /      Meeting     P|	�/V  �}	�/V  �m	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  �� /   �� /      Some_stuffs �	�/V  P�	�/V  ��	justforfun_justforfun_ 	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  Ю	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V  �uj /   �yj /      Appointment ��	�/V  0�	�/V  p�	Some_stuffs_Some_stuffs_ /V  ��	�/V  P�	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  0�	�/V  ��	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  �
�/V  �
�/V  ��	�/V  �	�/V  P 
�/V  �
�/V  
�/V  P
�/V  �
�/V  
�/V  �
�/V  

�/V  �
�/V  
�/V  �$
�/V  XԵ /   �Ե /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �� /   � /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               6�� /   ��� /       Meeting /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �h /   ��h /      Meeting     P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��� /    /      Workout     ��/V  p�/V  pThis_stuffs_This_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  j�� /   ��� /       Some_stuffs Ј�/V  P��/V  ЏSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  �, /   �, /   	   Meeting     ���/V  ���/V   �justforfun_justforfun_ �/V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  ��u /   �u /      Some_stuffs P�/V  ��/V  This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �o /   �o /      Meeting     �R�/V  �S�/V  UThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  썳 /   ��� /      Appointment ���/V  Д�/V  �justforfun_justforfun_ �/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  �� /   � /      Workout      ��/V  ���/V  ��justforfun_justforfun_ �/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  塗 /   ��� /      Meeting     �		�/V  �
	�/V  	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  ��X /   ��X /      Meeting     PZ	�/V  �[	�/V  `L	Some_stuffs_Some_stuffs_ /V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  .�f /   \�f /      Workout     ��	�/V  П	�/V  `�	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  Ю	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  \^x /   �^x /      Birthday V  �	�/V  0�	�/V  p�	This_stuffs_This_stuffs_ /V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  p�	�/V  @�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V   �	�/V  `�	�/V  ��	�/V  P�	�/V  ��	�/V  0�	�/V  p�	�/V  Q� /   �W� /       Meeting /V  P 
�/V  �
�/V  
This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  
�/V  �$
�/V  �%
�/V   
�/V  `
�/V  �
�/V  
�/V  P
�/V  �
�/V  P
�/V  �
�/V  �
�/V  
�/V  P
�/V  � 
�/V  "
�/V  :
�/V   '
�/V  `(
�/V  �)
�/V  �*
�/V   ,
�/V  �-
�/V   /
�/V  `0
�/V  �1
�/V  �f8 /   0g8 /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �+ /   ��* /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �� /   �� /      Appointment  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  1ou /   �pu /      Meeting     p��/V  ��/V  0�Some_stuffs_Some_stuffs_ /V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  p�/V  p�/V  DT� /   �X� /      Birthday    �#�/V  P%�/V  �)Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  Q� /   XR� /       Appointment ���/V   ��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  Ҳ� /   8�� /      Some_stuffs `��/V  ���/V  0�justforfun_justforfun_ �/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  q�Y /   (�Y /      Birthday    P�/V  ��/V  This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  $�K /   ��K /      Meeting     0H�/V  pI�/V  �JSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  0@� /   X@� /       Birthday    �~�/V   ��/V  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ��* /   ��* /       Workout     @��/V  ���/V  ��justforfun_justforfun_ �/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V  `� /   n� /      Workout     @��/V  � 	�/V  �	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  �Hw /   EEw /      Appointment @@	�/V  �A	�/V  �B	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  ؠK /   ڠK /      Birthday    �u	�/V  �v	�/V  `x	Some_stuffs_Some_stuffs_ /V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  �+ /   M+ /      Birthday    �	�/V  0�	�/V  p�	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  0�	�/V  p�	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  p�	�/V  @�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  r� /   � /      Meeting /V  ��	�/V  0�	�/V  p�	justforfun_justforfun_ 	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  �
�/V  �
�/V  ��	�/V  �	�/V  P 
�/V  �
�/V  
�/V  P
�/V  �
�/V  
�/V  �
�/V  

�/V  �
�/V  
�/V  �$
�/V  �%
�/V   
�/V  `
�/V  �
�/V  
�/V  P
�/V  �
�/V  P
�/V  5�� /   �� /      Some_stuffs "
�/V  :
�/V   '
Some_stuffs_Some_stuffs_ /V   ,
�/V  �-
�/V   /
�/V  `0
�/V  �1
�/V  `3
�/V  �4
�/V   6
�/V  �7
�/V  �N
�/V  P;
�/V  �<
�/V  >
�/V  �?
�/V  A
�/V  PB
�/V  �C
�/V  �D
�/V  F
�/V  PG
�/V  �H
�/V  �I
�/V  K
�/V  �L
�/V  �c
�/V  e
�/V  �O
�/V  0Q
�/V  pR
�/V  �W /   �W /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             E�w /   ,�w /      Workout /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �j� /   l� /      Workout     P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  J�� /   1�� /      Some_stuffs ��/V  p�/V  pThis_stuffs_This_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  Sٳ /   �ڳ /      Some_stuffs Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  �G- /   �B- /      Some_stuffs ���/V  ���/V   �Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  �+ /   ڙ+ /       Some_stuffs � �/V  0�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  �^< /   �f< /      Some_stuffs  <�/V  �F�/V  @?This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  n$� /   �)� /      Appointment 0s�/V  pt�/V  �uThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  �TK /   �XK /   	   Meeting     ���/V  Ъ�/V  P�justforfun_justforfun_ �/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V  �a� /   �a� /      Some_stuffs ���/V  ���/V  �Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  	"J /   �J /       Appointment @	�/V  �,	�/V  �	Some_stuffs_Some_stuffs_ /V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  �v /   �v /   	   Appointment �Q	�/V  �R	�/V  T	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  �+ /   ͼ+ /      Meeting     ��	�/V  Ж	�/V  �	Some_stuffs_Some_stuffs_ /V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  Ю	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  �� /   � /      Birthday V  ��	�/V   �	�/V  @�	Some_stuffs_Some_stuffs_ /V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V   �	�/V  `�	�/V  ��	�/V  P�	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  0�	�/V  ��	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  �
�/V  �
�/V  ��	�/V  �	�/V  P 
�/V  Q� /   V� /      Meeting /V  �
�/V  

�/V  �
justforfun_justforfun_ 
�/V   
�/V  `
�/V  �
�/V  
�/V  P
�/V  �
�/V  P
�/V  �
�/V  �
�/V  
�/V  P
�/V  � 
�/V  "
�/V  :
�/V   '
�/V  `(
�/V  �)
�/V  �*
�/V   ,
�/V  �-
�/V   /
�/V  `0
�/V  �1
�/V  `3
�/V  �4
�/V   6
�/V  �7
�/V  �N
�/V  P;
�/V  Z�� /   �� /      Workout /V  �C
�/V  �D
�/V  F
Some_stuffs_Some_stuffs_ /V  K
�/V  �L
�/V  �c
�/V  e
�/V  �O
�/V  0Q
�/V  pR
�/V  �S
�/V  �T
�/V  pV
�/V  �W
�/V  pY
�/V  �Z
�/V  0\
�/V  �]
�/V  0_
�/V  p`
�/V  �a
�/V  �z
�/V  �{
�/V  Pf
�/V  �g
�/V  i
�/V  Pj
�/V  �k
�/V  �l
�/V  n
�/V  Po
�/V  �p
�/V  �%) /   �%) /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             Tٳ /   0ڳ /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ��* /   Ы* /      Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ��g /   2�g /      Some_stuffs P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ,+; /   /+; /      Meeting     ��/V  p�/V  pjustforfun_justforfun_ �/V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  ţ9 /   ��9 /       Some_stuffs ���/V   ��/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  � X /   �X /      Appointment `��/V  ���/V  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  �� /   �� /       Workout     P�/V  ��/V  This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  ET� /   *X� /      Workout     0H�/V  pI�/V  �JSome_stuffs_Some_stuffs_ /V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �� /   � /      Appointment ���/V  0��/V  p�Some_stuffs_Some_stuffs_ /V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  �I /   =�I /      Birthday    ��/V  P��/V  ��justforfun_justforfun_ �/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  `�� /   :�� /      Meeting     �		�/V  �
	�/V  	justforfun_justforfun_ 	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  ��W /   Y�W /       Appointment @@	�/V  �A	�/V  �B	justforfun_justforfun_ 	�/V  �G	�/V  0I	�/V  PZ	�/V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  P�W /   �W /      Meeting     �u	�/V  �v	�/V  `x	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��	�/V   �	�/V  @�	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  YԵ /   �Ե /      Birthday    ��	�/V   �	�/V  p�	This_stuffs_This_stuffs_ /V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  p�	�/V  @�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��f /   �f /      Birthday     �	�/V  `�	�/V  ��	justforfun_justforfun_ 	�/V  p�	�/V  ��	�/V  0�	�/V  ��	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  �
�/V  �
�/V  ��	�/V  �	�/V  P 
�/V  �
�/V  
�/V  P
�/V  �
�/V  
�/V  �
�/V  

�/V  �
�/V  
�/V  �$
�/V  �%
�/V   
�/V  `
�/V  �
�/V  $�; /   ��; /      Some_stuffs �
�/V  
�/V  P
Some_stuffs_Some_stuffs_ /V   '
�/V  `(
�/V  �)
�/V  �*
�/V   ,
�/V  �-
�/V   /
�/V  `0
�/V  �1
�/V  `3
�/V  �4
�/V   6
�/V  �7
�/V  �N
�/V  P;
�/V  �<
�/V  >
�/V  �?
�/V  A
�/V  PB
�/V  �C
�/V  �D
�/V  F
�/V  PG
�/V  �H
�/V  �I
�/V  K
�/V  �L
�/V  �c
�/V  
 /   � /      Appointment �T
�/V  pV
�/V  �W
This_stuffs_This_stuffs_ /V  �]
�/V  0_
�/V  p`
�/V  �a
�/V  �z
�/V  �{
�/V  Pf
�/V  �g
�/V  i
�/V  Pj
�/V  �k
�/V  �l
�/V  n
�/V  Po
�/V  �p
�/V  Pr
�/V  �s
�/V  u
�/V  �v
�/V  �w
�/V  y
�/V  �
�/V  0}
�/V  p~
�/V  �
�/V  ��
�/V  0�
�/V  p�
�/V  ��
�/V  ?GZ /   MZ /      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     � /   � /      Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �Hw /   ,Kw /   	   Appointment  U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  i� /   F� /      Birthday    P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �%) /   �') /       Birthday    �#�/V  P%�/V  �)This_stuffs_This_stuffs_ /V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  �� /   �� /       Some_stuffs ���/V   ��/V  ��Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  � /   '� /      Meeting     `��/V  ���/V  0�This_stuffs_This_stuffs_ /V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  paW /   �aW /      Workout     �!�/V  #�/V  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V  ��u /   \�u /      Birthday    0]�/V  p^�/V  �_This_stuffs_This_stuffs_ /V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ��i /   �i /      Some_stuffs ���/V  Д�/V  �justforfun_justforfun_ �/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  �v /   �v /      Workout      ��/V  ���/V  ��This_stuffs_This_stuffs_ /V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  Xg /   �g /   	   Some_stuffs �		�/V  �
	�/V  	This_stuffs_This_stuffs_ /V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  �P� /   _J� /      Birthday    PZ	�/V  �[	�/V  `L	Some_stuffs_Some_stuffs_ /V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �I /   ��I /      Appointment ��	�/V  ��	�/V   �	Some_stuffs_Some_stuffs_ /V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  �1 /   �. /      Appointment �	�/V  0�	�/V  p�	Some_stuffs_Some_stuffs_ /V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  p�	�/V  @�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  � /   �� /      Birthday    ��	�/V  0�	�/V  p�	Some_stuffs_Some_stuffs_ /V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  �
�/V  �
�/V  ��	�/V  �	�/V  P 
�/V  �
�/V  
�/V  P
�/V  �
�/V  
�/V  �
�/V  

�/V  �
�/V  
�/V  �$
�/V  �%
�/V   
�/V  `
�/V  �
�/V  
�/V  P
�/V  �
�/V  P
�/V   8� /   "8� /      Birthday V  "
�/V  :
�/V   '
This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  `0
�/V  �1
�/V  `3
�/V  �4
�/V   6
�/V  �7
�/V  �N
�/V  P;
�/V  �<
�/V  >
�/V  �?
�/V  A
�/V  PB
�/V  �C
�/V  �D
�/V  F
�/V  PG
�/V  �H
�/V  �I
�/V  K
�/V  �L
�/V  �c
�/V  e
�/V  �O
�/V  0Q
�/V  pR
�/V  -+; /   �(; /      Appointment p`
�/V  �a
�/V  �z
justforfun_justforfun_ 
�/V  i
�/V  Pj
�/V  �k
�/V  �l
�/V  n
�/V  Po
�/V  �p
�/V  Pr
�/V  �s
�/V  u
�/V  �v
�/V  �w
�/V  y
�/V  �
�/V  0}
�/V  p~
�/V  �
�/V  ��
�/V  0�
�/V  p�
�/V  ��
�/V  ��
�/V  0�
�/V  ��
�/V  ��
�/V   �
�/V  ��
�/V   �
�/V  `�
�/V  D�� /   ^�� /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                      �: /   '�: /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     /�f /    �f /      Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �x /   �x /      Workout     ���/V  @��/V  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  �� /   �� /      Appointment �/�/V   1�/V  �5Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  P��/V  ���/V  `��/V   ��/V  �� /   ��� /      Some_stuffs ���/V   ��/V  @�This_stuffs_This_stuffs_ /V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  `��/V  0��/V  p��/V  ���/V  �� /   �� /      Meeting     ���/V  ���/V  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  ��, /   �, /      Birthday    ��/V  `�/V  �Some_stuffs_Some_stuffs_ /V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  퍳 /   #�� /      Workout     `M�/V  �N�/V  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ��w /   0�w /   	   Appointment ���/V  0��/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  �G- /   rK- /      Birthday     ��/V  `��/V  мSome_stuffs_Some_stuffs_ /V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  �[ /   ~[ /   	   Meeting     0��/V  ���/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V  ��h /   �h /      Appointment @3	�/V  �4	�/V  �5	Some_stuffs_Some_stuffs_ /V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �� /   �� /      Meeting     P|	�/V  �}	�/V  �m	Some_stuffs_Some_stuffs_ /V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  ��u /   ��u /      Meeting     ��	�/V  Щ	�/V  �	justforfun_justforfun_ 	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  P� /   z� /      Workout     p�	�/V  ��	�/V  ��	justforfun_justforfun_ 	�/V   �	�/V  `�	�/V  ��	�/V  P�	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  0�	�/V  ��	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  �
�/V  �
�/V  ��	�/V  �	�/V  P 
�/V  �
�/V  
�/V  P
�/V  �
�/V  
�/V  �
�/V  

�/V  �
�/V  "iJ /   poJ /      Appointment �
�/V  
�/V  P
justforfun_justforfun_ 
�/V  �
�/V  
�/V  P
�/V  � 
�/V  "
�/V  :
�/V   '
�/V  `(
�/V  �)
�/V  �*
�/V   ,
�/V  �-
�/V   /
�/V  `0
�/V  �1
�/V  `3
�/V  �4
�/V   6
�/V  �7
�/V  �N
�/V  P;
�/V  �<
�/V  >
�/V  �?
�/V  A
�/V  PB
�/V  �C
�/V  �D
�/V  F
�/V  �_� /   \_� /      Workout /V  �c
�/V  e
�/V  �O
This_stuffs_This_stuffs_ /V  �T
�/V  pV
�/V  �W
�/V  pY
�/V  �Z
�/V  0\
�/V  �]
�/V  0_
�/V  p`
�/V  �a
�/V  �z
�/V  �{
�/V  Pf
�/V  �g
�/V  i
�/V  Pj
�/V  �k
�/V  �l
�/V  n
�/V  Po
�/V  �p
�/V  Pr
�/V  �s
�/V  u
�/V  �v
�/V  �w
�/V  y
�/V  �
�/V  0}
�/V  ��� /   ߽� /   	   Birthday V  ��
�/V  ��
�/V  0�
This_stuffs_This_stuffs_ /V  ��
�/V   �
�/V  `�
�/V  ��
�/V  ��
�/V   �
�/V  P�
�/V  ��
�/V  Е
�/V  P�
�/V  ��
�/V  Й
�/V  �
�/V  ��
�/V  �
�/V  ��
�/V  Р
�/V  �
�/V  p�
�/V  ��
�/V  �
�/V  0�
�/V  @�
�/V  ��
�/V  @�
�/V  ��
�/V   �
�/V  @�
�/V  ��
�/V  �X /   ��X /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �G /   ��G /      Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �(� /   %� /      Meeting     P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �[ /   �	[ /   	   Some_stuffs ��/V  p�/V  pThis_stuffs_This_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  ��� /   J�� /   	   Meeting     Ј�/V  P��/V  ЏSome_stuffs_Some_stuffs_ /V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  �* /   �* /      Some_stuffs ���/V  ���/V   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  [' /   �& /      Birthday    `�/V  ��/V  �	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  p�V /   ��V /      Appointment @B�/V  �C�/V  PSome_stuffs_Some_stuffs_ /V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  桗 /   裗 /      Appointment �~�/V   ��/V  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  �+ /   � + /      Workout     ��/V  0��/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  �� /   � /      Birthday    ���/V   ��/V  @�This_stuffs_This_stuffs_ /V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V  