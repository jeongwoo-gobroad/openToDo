   
   ��7f    ˿7f    d       Test_Two                                P��U      Workout ffs  ��U  ���U  @ Some_stuffs_Some_stuffs_ �U  @"��U   #��U  �#��U  �$��U  ����U  P��U     Workout     ����U  @���U  �This_stuffs_This_stuffs_ �U  P���U  ���U   ���U  ����U  ����  us/       Birthday    @���U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  �9����  w/       Workout �U  ��	��U  P�	��U  ��	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �
��U  �g����  ��/      Appointment  o��U  �o��U  �pThis_stuffs_This_stuffs_ �U  Ps��U  t��U  �t��U  �u��U  ������  e�/       Meeting     ���U  `��U  Some_stuffs_Some_stuffs_ �U   ��U  ���U  ���U  ���U  �����  ��/       Birthday U  ����U  0���U  ��Some_stuffs_Some_stuffs_ �U  ����U  p���U  0���U  ����U  ����  ��/       Birthday    �n��U  po��U  0pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   t��U  �'����  Z�/      Meeting     ����U  @���U  ��Some_stuffs_Some_stuffs_ �U  ���U  @��U   ��U  ���U  ��S���  e/      Birthday nt �)��U  0*��U  �*This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p/��U  ������  �3/       Meeting      o��U  �o��U  �pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �u��U  $�����  84/      Appointment p���U  0���U  ��Some_stuffs_Some_stuffs_ �U  p��U  ���U  ���U  p��U  @�|���  h_/       Some_stuffs ����U  `���U  ��Some_stuffs_Some_stuffs_ �U  ���U  `��U  ��U  ���U  ����  �/       Appointment @.��U  �.��U  �/This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  �4��U  X&���  �/       Workout     ���U  0��U  �This_stuffs_This_stuffs_ �U  p��U  0��U  ���U  0��U  V�&���  ��/      Meeting     ����U  `���U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �c����  ��/       Meeting     ����U  p���U  0�Some_stuffs_Some_stuffs_ �U  ����U  0���U  ���U  ����U  �w����  ��/      Some_stuffs �/��U  p0��U  �4This_stuffs_This_stuffs_ �U  �>��U  �?��U   E��U  �F��U  �37���  ��/      Appointment ����U  ����U  @�Some_stuffs_Some_stuffs_ �U   ���U  ����U  0���U  ����U  �o����  -�/       Some_stuffs ����U  ����U  P�This_stuffs_This_stuffs_ �U  ���U  ����U  ����U  P���U  �����  �/      Some_stuffs p���U  ����U  ��This_stuffs_This_stuffs_ �U  0���U  ����U  ����U  0���U  pGe���  /       Birthday    ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  @���U  0���U   ���U  m3����  �&/      Birthday nt  ���U  ����U  @ This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  ����  5J/       Appointment Ю��U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  �I����  oo/       Meeting     ����U  P���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ����  $p/      Workout     p���U  ����U  ��This_stuffs_This_stuffs_ �U  p���U  ����U  p���U  ����U  ������  Nq/       Workout     ���U  ж��U  ��This_stuffs_This_stuffs_ �U  P���U  ���U  л��U  ����U  \�G���  ��/      Birthday    0A��U  �A��U  �BThis_stuffs_This_stuffs_ �U  0E��U  �E��U  pF��U  0G��U  �I����  H�/      Workout �U  p��U  0��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ������  +�/       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             Խi���  ��/      Meeting �U  0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  yw���  J�/       Meeting     ����U  @���U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `���U  �x���  !/       Some_stuffs Р��U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �����  4/      Meeting     ���U  ����U  P�Some_stuffs_Some_stuffs_ �U  @���U  ���U  ���U  ����U  +V���  �/       Some_stuffs  Q��U  �Q��U   RSome_stuffs_Some_stuffs_ �U  @T��U  �T��U  @U��U  �U��U  �����  �/       Workout     @S��U  �S��U  @TThis_stuffs_This_stuffs_ �U  @V��U   W��U  �W��U  @X��U  ����  _0/       Birthday    Т��U  P���U  �justforfun_justforfun_ ��U  Ц��U  ����U  ���U  Ш��U  \����  �0/      Appointment  ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  p���U  ���U  ж��U  �q����  �0/       Birthday    P���U  ���U  ��This_stuffs_This_stuffs_ �U  P���U  ����U  @��U  ���U  �7���  Z/       Workout �U  `���U   ���U  ��This_stuffs_This_stuffs_ �U  ����U  @���U   ���U  ����U  �1����  ��/       Birthday nt �|��U  p}��U  �}This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Ё��U  ������  �/      Appointment �Z��U  �[��U  @\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `a��U  J.i���  =�/       Workout     ����U  P���U  �Some_stuffs_Some_stuffs_ �U  P���U  ����U  ����U  P���U  �9k���  è/       Birthday nt `���U   ���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  ��y���  z�/      Workout     ����U  `���U   �Some_stuffs_Some_stuffs_ �U  `���U   ���U  ����U  ����U  :����  �/       Appointment  ���U  ����U   �justforfun_justforfun_ ��U  `���U  ���U  ����U  ���U  �	���  /�/      Some_stuffs 0f��U  �g��U  �iSome_stuffs_Some_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  1����  ^�/       Some_stuffs ����U  P���U  ��justforfun_justforfun_ ��U  ����U  P���U  ����U  ����U  x$����  ��/       Meeting     ����U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  zq����  �/       Meeting     P��U  ���U  PThis_stuffs_This_stuffs_ �U  ���U  �	��U  �"��U  p#��U  �Ч���  ��/       Some_stuffs л��U  ����U  ��justforfun_justforfun_ ��U  0���U  ���U  ����U  p���U  �.����  ��/      Meeting ffs ���U  ����U  �justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ����U  ��+���  �/      Meeting      ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��,���  �/       Birthday    @ ��U   ��U  �This_stuffs_This_stuffs_ �U  ��U  ���U  P��U  ���U  ��5���  $/       Birthday                       justforfun_justforfun_                                       3"6���  >/       Birthday    ����U  `���U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �%����  pF/       Birthday                       justforfun_justforfun_                                       ݣ����  [H/      Birthday     |��U  �|��U  �}Some_stuffs_Some_stuffs_ �U  `���U   ���U  ����U  `���U  I�Z���  i/       Appointment  V��U  �V��U  �WSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0[��U  ��j���  4m/      Workout      o��U  �o��U  �pSome_stuffs_Some_stuffs_ �U  Ps��U  t��U  �t��U  �u��U  H�����  ]�/       Some_stuffs                    Some_stuffs_Some_stuffs_                                     �����  c�/      Some_stuffs `���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  L����  A�/      Some_stuffs �t��U  �u��U  vThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `{��U  Qp$���  R�/       Appointment ���U  ����U  `�Some_stuffs_Some_stuffs_ �U  ����U  @���U   ���U  ����U  H55���  ��/       Workout �U  ��U  ���U  �justforfun_justforfun_ ��U  ���U  ���U  p��U  0��U  &:���  ��/      Some_stuffs ����U  ���U  ��justforfun_justforfun_ ��U   ���U  ����U  `���U  ����U  )"����  i/       Some_stuffs ���U  �	��U  �"Some_stuffs_Some_stuffs_ �U  ���U  p��U  0��U  ���U  d�����  @/      Birthday    p��U  0��U  0justforfun_justforfun_ ��U   +��U  �+��U  �/��U  p0��U  ������  �/       Workout     ����U  0���U  �This_stuffs_This_stuffs_ �U  0���U  ����U  0���U  ����U  �;s��  �#/       Meeting  U  ����U   ���U  ��justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ���U  �w��  !�#/       Appointment ����U  `���U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  H~��  յ#/       Meeting     �t��U  �u��U  vjustforfun_justforfun_ ��U  `y��U   z��U  �z��U  `{��U  �|��  $�#/       Meeting     ����U  ����U  �justforfun_justforfun_ ��U  ����U  ����U  @���U  ����U  �{���  ��#/       Appointment ���U  p��U  0Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ���U  <����  W�#/      Birthday U  Н��U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �#��  �#/       Meeting �U  @g��U  �g��U  �hjustforfun_justforfun_ _This_stuffs_This_stuffs_ �U   m��U  �Z*��  ��#/       Birthday nt 04��U  �4��U  05This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  p9��U  ̓-��  ��#/      Appointment ����U  @���U   �Some_stuffs_Some_stuffs_ �U  ���U  ж��U  ����U  P���U  |����  �$/      Workout     �*��U  P+��U  �+This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �/��U  \�;��  �'$/      Some_stuffs @���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��@��  #)$/       Some_stuffs `5��U  �5��U  `6This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ;��U  ��L��  C,$/       Meeting �U  �8��U  �9��U   :justforfun_justforfun_ ��U  0<��U  �<��U  0=��U  �=��U  qPR��  �-$/       Birthday    p��U  ���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p��U  �eU��  p.$/       Workout     @��U  ���U  ��Some_stuffs_Some_stuffs_ �U  p���U  ����U  p���U  ����U  4�W��  �.$/       Birthday    PF��U  �F��U  PGThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �K��U  �}���  �W$/      Some_stuffs ����U   ���U  ��justforfun_justforfun_ ��U  ����U  `���U  ���U  ����U  ��x��  y$/       Birthday    ���U  ����U  0�justforfun_justforfun_ ��U   ���U  ����U  ����U  @���U  �b���  $/      Meeting     0y��U  �y��U  pzjustforfun_justforfun_ ��U  �|��U  �}��U  0~��U  ����U  �
��  �$/      Some_stuffs @f��U  �f��U  @gThis_stuffs_This_stuffs_ �U  �i��U  @j��U   k��U  �k��U  Ø��  ��$/       Some_stuffs @��U  ���U  @Some_stuffs_Some_stuffs_ �U  @��U  ���U  @��U   ��U  !� ��  �$/       Meeting     ����U  0���U  �justforfun_justforfun_ ��U  0���U  ����U  0���U  ���U  �,!��  $�$/       Appointment �8��U  p9��U  �9This_stuffs_This_stuffs_ �U  P=��U  >��U  �>��U  ?��U  ����  9�$/       Some_stuffs                    This_stuffs_This_stuffs_                                     ����  ��$/       Appointment �U��U  �V��U  P[This_stuffs_This_stuffs_ �U  `f��U   g��U   l��U  �l��U  R�9 ��  ��$/       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             YBC ��  g�$/       Meeting     ����U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  p���U  0���U  ����U  �bJ ��  :�$/      Some_stuffs ���U  ����U  �justforfun_justforfun_ ��U  ����U  ���U  Ѕ��U  ����U  ��� ��  9%/       Meeting     ���U  @��U   This_stuffs_This_stuffs_ �U  0E��U  �E��U   ��U  ���U  ��� ��  :%/      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �T� ��  �%/       Appointment PC	��U  �C	��U  �D	Some_stuffs_Some_stuffs_ �U  �F	��U  PG	��U  �G	��U  �H	��U  q6h!��  f9%/       Workout     ����U  @���U  �Some_stuffs_Some_stuffs_ �U  P���U  ���U   ���U  ����U  �u!��  �<%/      Birthday    ����U  `���U  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  P�x!��  �=%/       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             r��!��  A%/       Some_stuffs �L��U  �M��U  @^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �R��U  ��"��  !h%/       Appointment  u��U  �u��U   vThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  z��U  d
�"��  @�%/      Appointment ����U   ���U  @�This_stuffs_This_stuffs_ �U  @���U   ���U  ����U  @���U  ���"��  Í%/       Meeting     �H��U  �I��U  0Jjustforfun_justforfun_ ��U  �L��U  �M��U  @^��U  �^��U  �=#��  ��%/      Appointment е��U  ����U  �Some_stuffs_Some_stuffs_ �U  ����U  ����U  ���U  ����U  �z�#��  <�%/      Meeting �U   �	��U  ��	��U   �	justforfun_justforfun_ 	��U   �	��U  ��	��U   �	��U  ��	��U  �8�#��  y�%/       Some_stuffs p���U  ����U  p�justforfun_justforfun_ ��U  ����U  p���U  0���U  ����U  �c$��  ��%/       Some_stuffs �m��U  @n��U  �nSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �s��U  S�k$��  ��%/       Birthday     g��U  �g��U   hSome_stuffs_Some_stuffs_ �U  �j��U  `k��U  �k��U  `l��U  ��q$��  � &/       Workout     ���U  ����U  P�Some_stuffs_Some_stuffs_ �U   ���U  ����U  P���U  ����U  ��$��  �&/      Workout     PH��U  I��U  �IThis_stuffs_This_stuffs_ �U  PL��U  M��U  �M��U  �N��U  `<
%��  |'&/       Workout     �G��U  0H��U  �Hjustforfun_justforfun_ ��U  �K��U  0L��U  �L��U  �M��U  ���%��  Q&/      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �?&��  �v&/      Some_stuffs �
��U  ���U  pThis_stuffs_This_stuffs_ �U  ���U  ���U  p��U  0��U  ��&��  ��&/       Appointment д��U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �f�&��  �&/       Meeting     �Y��U   Z��U  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @_��U  <�`'��  ��&/      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             y2|'��  ��&/       Birthday    �?��U  P@��U  AThis_stuffs_This_stuffs_ �U  �C��U  �D��U  E��U  �E��U  $	�'��  ��&/      Birthday     ���U  p���U  ��justforfun_justforfun_ ��U  ����U  `���U   ���U  ����U  �9�(��  q'/      Appointment ����U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  XG�(��  �'/       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ��(��  �'/       Some_stuffs ����U  `���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��1)��  �7'/      Workout     P[��U  \��U  �`This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �h��U  4,�)��  �^'/      Meeting      ���U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  P�a*��  ��'/       Some_stuffs ����U  @���U  �This_stuffs_This_stuffs_ �U  P���U  ���U   ���U  ����U  tci*��  ��'/       Workout �U  Я	��U  P�	��U  а	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��	��U  [�i*��  ��'/       Workout     p��U  ���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p$��U  2�o*��  �'/       Meeting ent ���U  P��U  �This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  p��U  M�r*��  �'/      Workout �U  ���U  ����U  @�This_stuffs_This_stuffs_ �U  p���U  ���U  ����U  P���U  �zx*��  c�'/       Some_stuffs �	��U  ��	��U  @�	Some_stuffs_Some_stuffs_ �U  p�	��U   �	��U  ��	��U   �	��U  ���*��  )�'/      Birthday     ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ж��U  @^�*��  h�'/       Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             4R�+��  B�'/      Appointment 0E��U  �E��U  pFSome_stuffs_Some_stuffs_ �U  �H��U  �I��U  0J��U  �J��U  i��+��  ��'/       Meeting ent �7��U   8��U  �_This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  0<��U  Y@W��  '�2/       Meeting ffs P���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��+W��  ��2/      Meeting     ����U  @���U  P�justforfun_justforfun_ ��U  P���U  Т��U  ����U  P���U  	p�W��  �3/       Birthday    ���U  0 ��U  � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0&��U  ظ�W��  w!3/       Some_stuffs �2��U   3��U   4Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `8��U  {3�W��  ["3/       Birthday    w��U  �w��U  xThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �|��U  B�W��  �$3/      Meeting     е��U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��CX��  �D3/      Birthday U  0���U  ����U  p�This_stuffs_This_stuffs_ �U  ����U   ���U  @���U   ���U  �KX��  �F3/       Birthday U   ���U  ����U  ��This_stuffs_This_stuffs_ �U  0���U  ����U  ����U  p���U  ��UX��  6I3/       Workout     ���U  ����U  `�Some_stuffs_Some_stuffs_ �U  ����U  `���U  ���U  ����U  8}�X��  �m3/       Some_stuffs @'��U  �'��U  @(This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �,��U  !b|Y��  ��3/       Meeting     ����U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  @���U   ���U  ����U  ���Y��  G�3/      Appointment �i��U  �j��U  `kSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   p��U  �q
Z��  �3/      Meeting     �Y��U   Z��U  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @_��U  �Z��  L�3/       Appointment ����U  `���U  ��Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  `���U  �,Z��  v�3/       Workout     @���U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  ��Z��  ��3/       Workout     ����U   ���U  ��justforfun_justforfun_ ��U  @���U  ����U  @���U  ����U  S�'Z��  r�3/       Meeting     ����U  @���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  .!�Z��  ��3/      Workout     ����U  p���U  0�justforfun_justforfun_ ��U  0���U  ����U  p���U  0���U  ��Z��  J�3/       Meeting                        justforfun_justforfun_ _                                     �l�Z��  v�3/       Some_stuffs �*��U  p+��U  0,This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �0��U  �K�Z��  ��3/       Meeting     `���U   ���U  ��Some_stuffs_Some_stuffs_ �U  `���U   ���U  ����U   ���U  �lB[��  �4/       Meeting     ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  �DH[��  O
4/       Some_stuffs ���U  `��U  �justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  �#��U  �'T[��  Z4/      Meeting     �|��U  �}��U  0~This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  l��[��  U34/      Some_stuffs �H��U  @I��U  �Ijustforfun_justforfun_ ��U  �K��U  @L��U  �L��U  �M��U  ��k\��  �T4/      Some_stuffs  E��U  �F��U  0KSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  \��U  ��n\��  �U4/       Meeting     ����U  P���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  [vs\��  �V4/       Some_stuffs ���U  p���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �|}\��  xY4/       Workout     �K��U  @L��U  �LThis_stuffs_This_stuffs_ �U  pO��U  �O��U  �P��U   Q��U  �]��  �{4/      Meeting     ���U  @	��U  �	Some_stuffs_Some_stuffs_ �U   ��U  ���U  @��U  ���U  8
]��  }4/       Meeting     ����U  `���U  ��justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ���U  �!]��  Y�4/       Appointment  -��U  �-��U   .Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   2��U  �¾]��  ��4/       Appointment  E��U  �F��U  0KThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  \��U  ��4^��  ��4/       Workout     ���U  ����U  `�justforfun_justforfun_ ��U  ����U  @���U   ���U  ����U  %�B^��  x�4/      Birthday    ���U  й��U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ���^��  ��4/      Some_stuffs                    Some_stuffs_Some_stuffs_                                     	��^��  ��4/       Workout      ���U  ����U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  ��i_��  5/       Workout     ���U  ����U  �Some_stuffs_Some_stuffs_ �U  Ѕ��U  ����U  ���U  ����U  $|�_��  �5/      Birthday    ����U  @���U  �This_stuffs_This_stuffs_ �U  P���U  ���U   ���U  ����U  J�_��  =?5/       Meeting ent  ���U  ����U  ��Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  �*`��  �A5/      Meeting �U  �}��U  ����U  pjustforfun_justforfun_ _ �U  p���U  0���U  ����U  ���U  �``��  yE5/       Appointment `���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  <)�`��  wg5/      Some_stuffs                    justforfun_justforfun_                                       �˱`��  m5/       Meeting ffs ����U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  ĽBa��  �5/      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             	rJa��  �5/       Some_stuffs `f��U   g��U   ljustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  �r��U  ��La��  ��5/       Appointment `/	��U  �/	��U  `0	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �3	��U  �V�a��  �5/       Workout     @���U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  ���a��  Q�5/      Appointment ���U  p��U  0Some_stuffs_Some_stuffs_ �U  �
��U  ���U  p��U  ���U  3�a��  �5/       Birthday nt �p��U  �q��U   rjustforfun_justforfun_ _ his_stuffs_This_stuffs_ �U  �u��U  {�a��  ��5/       Workout      E��U  �F��U  0KThis_stuffs_This_stuffs_ �U  �U��U  �V��U  P[��U  \��U  ��gb��  �5/      Workout �U  ����U  p���U  0�justforfun_justforfun_ ��U  ����U  ����U  p ��U  0��U  �c��  �6/       Meeting     Р��U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �lc��  S	6/      Appointment ����U  @���U  P�Some_stuffs_Some_stuffs_ �U  P���U  Т��U  ����U  P���U  ��c��  �-6/       Meeting ffs �6��U  P7��U  �7This_stuffs_This_stuffs_ �U   :��U  �:��U  0;��U  �;��U  Y�c��  �06/       Some_stuffs 0���U  ����U  �Some_stuffs_Some_stuffs_ �U  p���U  ����U  p���U  0���U  (�c��  �06/      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             e\.d��  �Q6/      Meeting     @���U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��;d��  �T6/       Birthday    ����U  ����U  @�Some_stuffs_Some_stuffs_ �U   ���U  ����U  ����U  @���U  ��Ld��  KY6/       Appointment 0U��U  �U��U  `Vjustforfun_justforfun_ ��U  @Y��U   Z��U  �Z��U  �[��U  ��d��  Zy6/       Workout      ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  `���U   ���U  ����U  0��d��  �z6/       Birthday                       This_stuffs_This_stuffs_                                     ���d��  $|6/       Appointment �{��U  0|��U  �|justforfun_justforfun_ ��U  `���U  ����U  `���U   ���U  %/�d��  �|6/      Birthday    p��U  0��U  �This_stuffs_This_stuffs_ �U  ���U  ���U  p��U  ���U  �]e��  .�6/      Some_stuffs ���U  ����U  �Some_stuffs_Some_stuffs_ �U  P���U  ����U  P���U  ����U  9^e��  J�6/       Birthday     >��U  �>��U  `?Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pC��U  yWde��  ۠6/       Birthday    ����U  0���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  af��  ��6/       Workout     p1��U  �1��U  �2This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �6��U  P>	f��  �6/       Appointment @(��U  �(��U  p)Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �-��U  ��f��  ��6/       Meeting     ����U  ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0���U  ��f��  9�6/       Birthday    0��U  ���U  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  |�Ag��  7/      Meeting     E��U  �E��U  PFThis_stuffs_This_stuffs_ �U  PH��U  I��U  �I��U  �J��U  �]h��  �c7/      Some_stuffs ���U  ����U  0�This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  @���U  �'eh��  �e7/       Some_stuffs P���U  ����U  P�Some_stuffs_Some_stuffs_ �U  ����U  p���U  ����U  p���U  :xqh��  �h7/       Birthday    k	��U  �k	��U  l	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �o	��U  ��h��  <�7/      Meeting     P���U  ���U  Цjustforfun_justforfun_ ��U  ����U  P���U  Ъ��U  ����U  ��i��  �7/       Appointment                    justforfun_justforfun_                                        l����  �;B/       Birthday    0���U  ����U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  vA���  �^B/       Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �I���  �`B/      Some_stuffs ����U  `���U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �CL���  YaB/       Appointment @\��U  �\��U  @]This_stuffs_This_stuffs_ �U  �_��U  �`��U   a��U  �a��U  �+ܓ��  0�B/      Birthday U  0f��U  �g��U  �iSome_stuffs_Some_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  �����  .�B/       Some_stuffs `V��U   W��U  �WThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ]��U  6�p���  B�B/      Some_stuffs 0�	��U  ��	��U  0�	Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ��	��U  q�p���  F�B/       Appointment b��U  �b��U  PcThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �g��U  ��x���  6�B/       Some_stuffs ����U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  k���  ��B/      Appointment ���U  ����U  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �w���  /�B/       Appointment �t��U  �u��U  vjustforfun_justforfun_ ��U  `y��U   z��U  �z��U  `{��U  f����  `�B/      Workout �U  ���U  ����U  p�This_stuffs_This_stuffs_ �U  ����U  P���U  ����U  P���U  �\����  ��B/       Meeting     ����U  ����U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  �����  C C/       Appointment �<��U  �=��U   >This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �A��U  2Q;���  �!C/       Some_stuffs 0��U  ���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �$��U  �<���  
"C/       Appointment pF��U  0G��U  �Gjustforfun_justforfun_ ��U  0J��U  �J��U  �K��U  0L��U  �xD���  �#C/       Some_stuffs p���U  ���U  ��This_stuffs_This_stuffs_ �U  0���U  ����U  ����U  0���U  �K���  �%C/       Birthday U  ����U  ����U  �Some_stuffs_Some_stuffs_ �U  ���U  ����U  P���U  ����U  � X���  �(C/       Birthday     ���U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  �]���  l*C/       Appointment  ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ����  pLC/      Birthday nt �z��U  `{��U   |This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  �o���  hpC/      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �;���  ,�C/       Workout     ����U  p���U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0��U  �!���  .�C/      Birthday    `���U   ���U  ��Some_stuffs_Some_stuffs_ �U   ���U  ����U  `���U   ���U  ������  n�C/       Meeting     p?��U  �?��U  p@justforfun_justforfun_ ��U  �B��U  pC��U  �C��U  �D��U  �ɲ���  F�C/      Meeting     Н��U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  Ȣ����  �C/       Workout     `_��U   `��U  �`Some_stuffs_Some_stuffs_ �U   c��U  �c��U  `d��U  �d��U  B�=���  ��C/       Meeting ffs  f��U  �f��U   gThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  `k��U  �YN���  �C/       Some_stuffs  +��U  �+��U  �/This_stuffs_This_stuffs_ �U  �9��U  �:��U  �>��U  �?��U  �hT���  ��C/      Appointment �B��U  PC��U  �Cjustforfun_justforfun_ ��U  PF��U  �F��U  PG��U  �G��U  )hV���  )�C/       Birthday    ���U  0��U  �This_stuffs_This_stuffs_ �U  p��U  0��U  ���U  0��U  �����  �D/       Meeting �U  ����U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  u����  *D/      Workout     �t��U  �u��U  vThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `{��U  ����  �D/       Workout ent P���U  ���U  лSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �w���  D7D/      Meeting     ���U  ����U  P�This_stuffs_This_stuffs_ �U  @���U  ���U  ���U  ����U  ��}���  �8D/       Workout     �w��U  px��U  0ySome_stuffs_Some_stuffs_ �U  �{��U  0|��U  �|��U  �}��U  :�����  �;D/       Meeting     pv��U  0w��U  �wThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0|��U  �L#���  &cD/      Meeting     �R��U  PS��U  TSome_stuffs_Some_stuffs_ �U  �q��U  `r��U   W��U  �W��U  1�����  ��D/       Some_stuffs ����U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  <S����  ��D/      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �=����  A�D/       Workout �U  0���U  ���U  ��Some_stuffs_Some_stuffs_ �U  ���U  p���U  0���U  ����U  y7���  ۩D/       Birthday U  0f��U  �g��U  �iSome_stuffs_Some_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  �K���  ܮD/      Some_stuffs �g��U  �h��U  pjThis_stuffs_This_stuffs_ �U  �m��U  @n��U   o��U  �o��U  $�ܜ��  8�D/      Some_stuffs Ц��U  ����U  �This_stuffs_This_stuffs_ �U  Ъ��U  ����U  P���U  ���U  �Ip���  ��D/       Workout     ����U  ����U  p�Some_stuffs_Some_stuffs_ �U  0���U  ����U  0���U  ����U  eZy���  @�D/      Meeting     �t��U  �u��U  vSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `{��U  XȀ���  '�D/       Meeting     ����U  ����U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  `���  �#E/       Meeting     �,��U  �-��U  @.This_stuffs_This_stuffs_ �U   1��U  �1��U  �2��U   3��U  򳜞��  �FE/       Meeting     л��U  ����U  ��justforfun_justforfun_ ��U  0���U  ���U  ����U  p���U  ������  �GE/      Appointment �z��U  `{��U   |justforfun_justforfun_ ��U  p��U  0���U  ����U  ����U  �ӥ���  ,IE/       Meeting     ����U  @���U  ��This_stuffs_This_stuffs_ �U  ���U  й��U  p���U  0���U  �ǩ���  /JE/       Meeting �U  ���U  p��U  0justforfun_justforfun_ ��U  ���U  0 ��U  � ��U  �!��U  �SI���  sE/      Some_stuffs ����U  @���U  �This_stuffs_This_stuffs_ �U  P���U  ���U   ���U  ����U  ��K���  �sE/       Some_stuffs p���U  ����U  ��justforfun_justforfun_ ��U  0���U  ����U  ����U  0���U  �#O���  �tE/       Workout                        This_stuffs_This_stuffs_                                     �ҟ��  *�E/       Appointment ����U  p���U  0�This_stuffs_This_stuffs_ �U  ���U  p���U  ���U  p���U  0�؟��  ��E/       Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �Oޟ��  +�E/       Some_stuffs ����U  `���U  ��Some_stuffs_Some_stuffs_ �U  0���U  ����U  p���U  ����U  �3���  0�E/      Birthday    �-	��U   .	��U  �q	Some_stuffs_Some_stuffs_ �U  `0	��U  �0	��U  `1	��U  �1	��U  b�^���  ��E/       Workout     `���U  ����U  `�justforfun_justforfun_ ��U  ����U   ���U  ����U  `���U  \Wl���  ��E/       Birthday    ���U  ����U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  Q�p���  ��E/       Meeting     ����U  `���U  ��This_stuffs_This_stuffs_ �U  `���U  ���U  ����U  ���U  �~���  D�E/      Workout     ����U  @���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  c����  |�E/       Meeting     �g��U  �h��U  pjThis_stuffs_This_stuffs_ �U  �m��U  @n��U   o��U  �o��U  rd����  &�E/       Some_stuffs ����U  @���U  ЋThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  v	���  ��E/       Some_stuffs �}��U  ����U  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  �����  ��E/       Some_stuffs                    justforfun_justforfun_                                       ����  ��E/      Some_stuffs ����U  @���U  P�Some_stuffs_Some_stuffs_ �U  P���U  Т��U  ����U  P���U  �#0���  01F/       Some_stuffs �Y��U   Z��U  �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @_��U  Ξ1���  �1F/      Workout ffs �o��U   p��U  �pThis_stuffs_This_stuffs_ �U   s��U  �s��U   t��U  �t��U  � D���  N6F/       Birthday    ����U  ���U  Тjustforfun_justforfun_ ��U  P���U  ���U  Ц��U  ����U  o����  �UF/       Meeting     ���U  0��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0��U  T�Ţ��  rWF/       Workout     ����U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @��U  "�ˢ��  YF/       Meeting     05��U  �5��U  06This_stuffs_This_stuffs_ �U  �8��U  p9��U  �9��U  �:��U  =�֢��  �[F/      Some_stuffs 0f��U  �g��U  �iSome_stuffs_Some_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  �ߢ��  ^F/       Meeting     �f��U  �g��U  `hSome_stuffs_Some_stuffs_ �U  `k��U   l��U  �l��U  `m��U  1^���  ~~F/       Some_stuffs P���U  ���U  ��justforfun_justforfun_ ��U  ����U  ����U  ���U  ����U  0�z���  ޅF/       Some_stuffs p��U  0��U  0This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p0��U  ������  ץF/       Workout     �N��U  PO��U  0Ajustforfun_justforfun_ ��U  0D��U  �D��U  0E��U  �E��U  �>����  ��F/       Appointment �<��U  �=��U   >Some_stuffs_Some_stuffs_ �U  �N��U  PO��U  0A��U  �A��U  46���  ¨F/      Workout ent                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             S���  �F/       Meeting     Ѕ��U  ����U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  Ћ��U  �+K���  �{Q/      Meeting     0y��U  �y��U  pzjustforfun_justforfun_ ��U  �|��U  �}��U  0~��U  ����U  ������  Y�Q/       Some_stuffs ���U  Ѓ��U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  Ј��U  \ku���  �Q/      Birthday U  0f��U  �g��U  �iSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �t��U  B����  ��Q/       Appointment 0���U  ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  )	����  ��Q/       Birthday U  0��U  ���U  �Some_stuffs_Some_stuffs_ �U  0��U  ���U  p��U  0��U  �<���  ~�Q/      Meeting                        justforfun_justforfun_                                       k���  ��Q/       Workout     p��U  0��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p��U  �$���  ��Q/       Birthday fs 0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  (�*���  i�Q/       Birthday nt P���U  ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  ������  DR/       Appointment                    Some_stuffs_Some_stuffs_                                     %����  xR/      Appointment p��U  0��U  0This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p0��U  �����  �hR/      Birthday    ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  ������  lR/       Meeting �U  0��U  ���U  �This_stuffs_This_stuffs_ �U  0��U  ���U  p��U  0��U  �x���  Q�R/      Appointment �|��U  �}��U  0~This_stuffs_This_stuffs_ �U  `���U   ���U  ����U  `���U  ����  ��R/      Some_stuffs                    justforfun_justforfun_                                       de����   �R/      Appointment 0���U   ���U  @�This_stuffs_This_stuffs_ �U  p���U  0���U  ����U  `���U  ��<���  .S/       Some_stuffs ���U  p��U  0justforfun_justforfun_ ��U  ���U  p��U  0��U  ���U  ��<���  ;S/      Meeting �U  �|��U  �}��U  0~Some_stuffs_Some_stuffs_ �U  `���U   ���U  ����U  `���U  TS���  �S/       Meeting      ���U  ����U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  H�����  )S/       Meeting     ����U  p���U  0�justforfun_justforfun_ ��U  ���U  ����U  ����U  @���U  �U����  �.S/      Appointment p��U  ���U  �This_stuffs_This_stuffs_ �U  ���U  @��U   ��U  ���U  �����  �/S/       Some_stuffs P���U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  ��u���  [QS/      Birthday     ���U  ����U  ��justforfun_justforfun_ ��U  ����U  p���U  ���U  ж��U  2}���  @SS/       Appointment  3��U  �3��U   4This_stuffs_This_stuffs_ �U  �6��U   7��U  �7��U   8��U  ",���  �vS/       Some_stuffs ����U  ���U  Тjustforfun_justforfun_ ��U  P���U  ���U  Ц��U  ����U  !���  xS/       Birthday    ����U  @���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �l#���  �}S/       Meeting     @���U    ��U  �This_stuffs_This_stuffs_ �U  ���U  P��U   ��U  ���U  tQ%���  J~S/      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ԡ���  *�S/       Workout     ����U  ����U   �justforfun_justforfun_ ��U  Ћ��U  ����U   ���U  ����U  �����  ��S/       Appointment 0D��U  �D��U  0ESome_stuffs_Some_stuffs_ �U  �G��U  0H��U  �H��U  �I��U  $����  ��S/       Appointment ����U  P���U  �justforfun_justforfun_ ��U  ����U  `���U  Э��U  P���U  6C����  �S/      Appointment  ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  hk����  ��S/       Birthday U  0f��U  �g��U  �iSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �t��U  j�8���  ��S/       Birthday fs 0�	��U  ��	��U  ��	Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  Њ	��U  6;���  n�S/      Meeting     p��U  0��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ��T���  ��S/       Some_stuffs ����U  P���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ������  ��S/       Some_stuffs �9��U  �:��U  �>Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @Q��U  �����  ��S/      Some_stuffs �[��U  `\��U  �\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @a��U  �\|���  �T/       Birthday    p���U  0���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  �����  (?T/      Meeting      ���U  ����U  �rThis_stuffs_This_stuffs_ �U  �u��U  v��U  �v��U  �w��U  �K����  �dT/       Birthday    '	��U  �'	��U  (	This_stuffs_This_stuffs_ �U  �*	��U   +	��U  �+	��U   ,	��U  �eL���  p�T/       Appointment                    justforfun_justforfun_                                       x����  ۭT/       Appointment `���U  �.	��U  `�justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ���U  ��l���  E�T/      Some_stuffs ���U  0��U  �This_stuffs_This_stuffs_ �U  ���U  ���U  p��U  0��U  �.q���  d�T/       Appointment @��U  ���U  @justforfun_justforfun_ _ �U  `��U   ��U  ���U   ��U  �\w���  ��T/       Meeting  fs 0��U  ���U  �This_stuffs_This_stuffs_ �U  0��U  ���U  ���U  0 ��U  ������  C#U/       Birthday    p��U  0��U  0This_stuffs_This_stuffs_ �U   +��U  �+��U  �/��U  p0��U  ������  �'U/      Appointment �z��U  `{��U   |justforfun_justforfun_ ��U  p��U  0���U  ����U  ����U  �-���  %KU/      Meeting     ����U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �3���  �LU/       Some_stuffs `f��U   g��U   lThis_stuffs_This_stuffs_ �U  pj��U  0k��U  �q��U  �r��U  ������  �xU/       Workout     ����U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  p���U  0���U  ����U  H����  �xU/       Workout      V��U  �V��U  �WSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0[��U  �c���  �U/       Some_stuffs ���U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �]{���  ��U/      Birthday    ����U  P���U  �justforfun_justforfun_ ��U  P���U  ����U  ����U  P���U  �����  )�U/      Meeting     ���U  0 ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �3��U  ]����  +�U/      Workout     �t��U  �u��U  vjustforfun_justforfun_ ��U  `y��U   z��U  �z��U  `{��U  ������  0�U/       Some_stuffs 05��U  �5��U  06Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �:��U  �v<���  �V/      Appointment  ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  )G���  IV/       Appointment �g��U  �h��U  pjThis_stuffs_This_stuffs_ �U  �m��U  @n��U   o��U  �o��U  D��	��  l�`/      Appointment                    justforfun_justforfun_                                       M}
��  ��`/      Appointment P���U  ���U  ��justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  @���U  �h~
��  ��`/       Birthday    0(��U  �(��U  �)justforfun_justforfun_ ��U  0,��U  �,��U  p-��U  0.��U  ���
��  ��`/       Some_stuffs ��	��U   �	��U  ��	This_stuffs_This_stuffs_ �U  ��	��U  `�	��U  �	��U  ��	��U  �,��  �a/      Birthday U  ����U  P���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��,��  �a/       Meeting     �g��U  �h��U  pjjustforfun_justforfun_ ��U  �m��U  @n��U   o��U  �o��U  �����  /5a/       Appointment `k��U   l��U  �lThis_stuffs_This_stuffs_ �U  `o��U   p��U  �p��U  �q��U  ����  :5a/       Some_stuffs ����U  ����U  `�justforfun_justforfun_ ��U   ���U  ���U  ����U  ���U  3Y���  �6a/       Meeting     ����U  `���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �����  �7a/       Meeting �U  �z��U  `{��U   |Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ����  �9a/       Birthday                       Some_stuffs_Some_stuffs_                                     9R��  �\a/       Meeting     �/��U  p0��U  �4justforfun_justforfun_ ��U  �>��U  �?��U   E��U  �F��U  ,�_��  -`a/      Some_stuffs ����U  @���U  P�Some_stuffs_Some_stuffs_ �U  P���U  Т��U  ����U  P���U  HM���  ��a/       Workout     PJ	��U  �J	��U  PK	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  O	��U  �s���  ��a/      Birthday fs ��	��U  `�	��U  ��	Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  `�	��U  ����  �a/      Workout     ���U   ��U  �justforfun_justforfun_ ��U   ��U  ���U   ��U  ���U  m���  �a/      Meeting     ����U  P���U  �justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  P���U  ��!��  Y�a/       Appointment  E��U  �F��U  0Kjustforfun_justforfun_ ��U  �U��U  �V��U  P[��U  \��U  |z���  ��a/      Birthday    ����U  `���U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  I����  ��a/       Meeting     `���U   ���U  ��justforfun_justforfun_ ��U   ���U  ����U  `���U   ���U  �*B��  :b/       Birthday    ����U  P���U  �This_stuffs_This_stuffs_ �U  ����U  P���U   ���U  ����U  �L��  �b/       Birthday    ����U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  ,	T��  �!b/      Appointment ���U  ����U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  :W��  �"b/       Birthday    ����U  `���U   �justforfun_justforfun_ _ �U  ����U  p���U  0���U  ����U  y!Y��  #b/       Appointment ����U  @���U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  �r��  kb/       Appointment @p��U   q��U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  v��U  \u���  Krb/      Meeting ffs ���U  P��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p��U  �w"��  /�b/       Workout ent �Y��U  0Z��U  �ZThis_stuffs_This_stuffs_ �U  �\��U  `]��U  ^��U  �^��U  `���  \�b/       Some_stuffs 0���U  ����U  p�justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U   ���U  #[���  4�b/       Birthday    ����U  ���U  ��Some_stuffs_Some_stuffs_ �U  @���U   ���U  ����U  @���U  Y����  '�b/       Some_stuffs �l��U  `m��U   This_stuffs_This_stuffs_ �U  �p��U  �q��U  0r��U  �r��U  D����  (�b/       Appointment �|��U  p}��U  �}justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  Ё��U  np���  վb/      Some_stuffs ����U  0���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  :��  ��b/       Meeting     ����U   ���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  !�<��  t�b/       Workout     �2��U   3��U   4Some_stuffs_Some_stuffs_ �U  `6��U   7��U  �7��U  `8��U  ��<��  ��b/       Appointment ����U  P���U   �justforfun_justforfun_ _ �U  @��U  ���U  ����U  0���U  ��G��  M�b/       Workout     P���U  ���U  РThis_stuffs_This_stuffs_ �U  ����U  P���U  ���U  ����U  
'���  5c/       Appointment ����U  @���U  �This_stuffs_This_stuffs_ �U  P���U  ���U   ���U  ����U  ty���  Jc/      Workout �U  0���U   ���U  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `���U  �����  �	c/       Meeting ent px��U  �x��U  pySome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p}��U  �����  �
c/       Appointment  o��U  �o��U  �pSome_stuffs_Some_stuffs_ �U  Ps��U  t��U  �t��U  �u��U  ��r��  �/c/       Workout                        This_stuffs_This_stuffs_                                     �nt��  =0c/      Birthday    ����U  `���U  ��justforfun_justforfun_ ��U  ���U  `��U  ��U  ���U  ����  95c/       Meeting      ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  `���U  ����U  `���U  4���  �[c/      Appointment p���U  0���U  ��justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  P���U  �P���  �~c/       Appointment p��U  0��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  d�B��  ��c/      Meeting     ����U  `���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  BG��  ��c/       Meeting      ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  �����  �c/       Appointment Т��U  P���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Ш��U   ����  ��c/       Appointment                    justforfun_justforfun_                                       �����  ��c/       Workout     ���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  �d��  ��c/      Some_stuffs 0���U   ���U  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `���U  �.��  �d/      Birthday    @���U   ���U  ��This_stuffs_This_stuffs_ �U  ����U  @���U   ���U  ����U  ���  yd/       Workout     ����U  0���U  ��justforfun_justforfun_ ��U  0���U  ����U  p���U  0���U  �z���  >Ed/      Workout �U  е��U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �F���  7Fd/       Birthday    �w��U  �x��U  PsSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �~��U  ����  nFd/       Meeting     0���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  v.��  �ed/      Some_stuffs `���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ��5��  �gd/       Appointment е��U  ����U  �This_stuffs_This_stuffs_ �U  ����U  ����U  ���U  ����U  �>M��  �md/       Meeting ffs ����U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  ����U  @���U   ���U  �����  ��d/      Birthday    ����U  `���U  ��This_stuffs_This_stuffs_ �U  ���U  `��U  ��U  ���U  �+���  ,�d/       Workout     �g��U  �h��U  pjjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  �o��U  �d��  C�d/       Meeting      ���U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  �nw��  9�d/       Meeting     ����U  p���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  9���  ��d/       Meeting     �C��U  �D��U  @EThis_stuffs_This_stuffs_ �U  �G��U   H��U  �H��U  @I��U  8���  ��d/       Appointment ���U   ��U  �Some_stuffs_Some_stuffs_ �U   ��U  ���U  0��U  ���U  �_���  �e/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ����  te/      Meeting ent ���U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  �,��  %*e/      Birthday    ����U  @���U  Ћjustforfun_justforfun_ ��U  ����U  `���U   ���U  ����U  U�wE��  ��o/      Workout �U  @���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  B�zE��  ��o/       Meeting     ����U   ���U  ��This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U   ���U   ��E��   p/       Some_stuffs 0f��U  �g��U  �iSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �t��U  �dF��  z%p/       Meeting     PO��U  �O��U  �PSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  �T��U  @5#F��  �)p/       Birthday                       Some_stuffs_Some_stuffs_                                     ��(F��  A+p/       Some_stuffs 0J��U  �J��U  �Kjustforfun_justforfun_ _ �U  @^��U  �^��U  �O��U  pP��U  �1F��  �-p/       Meeting     @���U  ����U  @�This_stuffs_This_stuffs_ �U  ����U   ���U  ����U  ����U  m2F��  �-p/      Appointment `f��U   g��U   lThis_stuffs_This_stuffs_ �U  pj��U  0k��U  �q��U  �r��U  h��F��  QPp/       Some_stuffs ����U  @���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ~�F��  �Pp/      Some_stuffs ����U  @���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0���U  � ]G��  %zp/      Appointment  ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  �R�G��  >�p/      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             *e�G��  I�p/       Workout     p���U  ���U  p�justforfun_justforfun_ ��U  ����U  0���U  ���U  ����U  ��G��  ˠp/       Workout     �<��U  �=��U   >Some_stuffs_Some_stuffs_ �U  �N��U  PO��U  0A��U  �A��U  ��{H��  ��p/      Meeting     ����U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  aI��  ��p/       Appointment �N��U  PO��U  0ASome_stuffs_Some_stuffs_ �U  0D��U  �D��U  0E��U  �E��U  �I��  T�p/      Some_stuffs �}��U  ����U  pSome_stuffs_Some_stuffs_ �U  p���U  0���U  ����U  ���U   �&I��  T�p/       Birthday    ����U  @���U  ��Some_stuffs_Some_stuffs_ �U  ����U  @���U  Ћ��U  ����U  �#.I��  0�p/       Birthday    �}��U  `~��U   This_stuffs_This_stuffs_ �U  ����U  `���U  ����U  `���U  r�I��  Dq/      Workout      ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  `���U   ���U  ����U  ���I��  �q/       Birthday    P���U  ���U  ��justforfun_justforfun_ ��U  ���U  ����U  P���U  ���U  `'�I��  \q/       Workout                        justforfun_justforfun_                                       �SJ��  L<q/       Meeting     ����U  @���U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  ��SJ��  O<q/       Appointment ����U   ���U  ��justforfun_justforfun_ ��U  ����U  `���U   ���U  ���U  !�SJ��  T<q/       Some_stuffs 0r��U  �r��U  �sThis_stuffs_This_stuffs_ �U  pv��U  0w��U  �w��U  px��U  ��XJ��  �=q/      Some_stuffs ����U  @���U  �This_stuffs_This_stuffs_ �U  P���U  ���U   ���U  ����U  "`_J��  T?q/       Appointment �t��U  Pu��U  �uSome_stuffs_Some_stuffs_ �U  x��U  �x��U  �y��U   z��U  ���J��  +_q/       Appointment 0��U  ���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0 ��U  ���J��  (`q/      Appointment ����U  `���U   �Some_stuffs_Some_stuffs_ �U  `���U  ����U  ����U  p���U  x��J��  {aq/       Birthday U  ���U  ж��U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ���K��  Z�q/       Some_stuffs ����U  `���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ��K��  j�q/       Birthday U  `���U   ���U  ��This_stuffs_This_stuffs_ �U  `���U   ���U  ����U  `���U  �x�K��  ��q/       Workout                        Some_stuffs_Some_stuffs_                                     `YL��  ��q/       Some_stuffs @���U    ��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  QCL��  2�q/       Some_stuffs p��U  0��U  �This_stuffs_This_stuffs_ �U  ���U  ���U  p��U  ���U  .�!L��  ��q/      Meeting      ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  ���L��  ��q/      Appointment                    justforfun_justforfun_                                       (a�L��  ��q/       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             l�L��  ��q/       Some_stuffs ���U  ����U  0�This_stuffs_This_stuffs_ �U   ���U  ����U  ����U  @���U  #[�L��  4�q/       Birthday    E��U  �E��U  PFSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �J��U  ���L��  b�q/       Workout      E��U  �F��U  0KThis_stuffs_This_stuffs_ �U  �U��U  �V��U  P[��U  \��U  )SHM��  	�q/       Some_stuffs �L��U  �M��U  @NThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   R��U  <JM��  w�q/      Birthday nt м��U  P���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  t��M��  
#r/      Some_stuffs p��U  0��U  0justforfun_justforfun_ ��U   +��U  �+��U  �/��U  p0��U  2-�M��  #r/       Birthday U  ����U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ���M��  �%r/       Appointment `6��U   7��U  �7Some_stuffs_Some_stuffs_ �U  `:��U   ;��U  �;��U  `<��U  9jN��  3Hr/       Some_stuffs �t��U  �u��U  vThis_stuffs_This_stuffs_ �U  `y��U   z��U  �z��U  `{��U  ��wN��  �Kr/      Workout     ����U  ����U  p justforfun_justforfun_ ��U  ���U  p��U  0��U  ���U  �~O��  rr/       Meeting     p���U  0���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  ��O��  $sr/       Meeting     p��U  ���U  �justforfun_justforfun_ ��U  p��U  0��U  ���U  ���U  �O��  ��r/       Some_stuffs @Y��U   Z��U  �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   `��U  ql�O��  &�r/       Meeting �U  0f��U  �g��U  �iThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �t��U  ��O��  %�r/       Workout                        Some_stuffs_Some_stuffs_                                     �?�O��  ��r/      Workout     ����U  `���U  @�justforfun_justforfun_ ��U  ����U  ����U  ����U  `���U  y�2P��  �r/       Appointment P���U  ���U  иSome_stuffs_Some_stuffs_ �U  ����U  P���U  м��U  P���U  �BP��  C�r/      Some_stuffs �Y��U   Z��U  �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @_��U  e�P��  ��r/       Some_stuffs 0���U  ����U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  �?�P��  Z�r/      Some_stuffs �t��U  �u��U  vSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `{��U  �Q��  �s/       Meeting      E��U  �F��U  0KThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  \��U  �^�Q��  s/       Appointment @���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  ��R��  �6s/       Some_stuffs p���U  ���U  ��This_stuffs_This_stuffs_ �U  0���U  ����U  ����U  0���U  %�R��  87s/      Meeting �U   V��U  �V��U  �Wjustforfun_justforfun_ ��U  �Y��U  0Z��U  �Z��U  0[��U  �R��  d\s/      Some_stuffs pR��U  �R��U  �SThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �X��U  �MS��  z�s/       Workout     ����U  @���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  k�S��  ��s/      Appointment p)��U  *��U  �*Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @/��U  ��S��  l�s/       Meeting     �c��U  �d��U  0eSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pj��U  �$rT��  ~�s/      Appointment ����U  ����U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �$	U��  &�s/      Appointment  ���U  ����U  `�justforfun_justforfun_ _ �U  ����U  ����U  `���U  ����U  H��U��  ]t/       Workout     @.��U  �.��U  �/Some_stuffs_Some_stuffs_ �U  �2��U   3��U   4��U  �4��U  t��U��  & t/       Birthday     E��U  �F��U  0KSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  \��U  ���U��  E!t/       Meeting     ����U  p���U  �Some_stuffs_Some_stuffs_ �U  @���U  ����U  @���U  ���U  ��U��  �$t/      Appointment �r��U  �s��U  @tjustforfun_justforfun_ _This_stuffs_This_stuffs_ �U  �x��U  !ܯU��  �$t/       Workout ffs �T��U  `U��U   VThis_stuffs_This_stuffs_ �U  �X��U  Y��U  �Y��U  0Z��U  ��,V��  �Dt/      Some_stuffs �i��U  �j��U  `kSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U   p��U  9�CV��  �Jt/       Some_stuffs P���U  ���U  ��Some_stuffs_Some_stuffs_ �U  ���U  о��U  ����U  P���U  ȕHV��  �Kt/       Meeting     ����U  ����U  P�justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ���U  �KV��  �Lt/       Appointment ����U  ���U  ��This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ���U  ��V��  Znt/      Workout     ����U  ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  ���V��  pt/       Appointment � ��U  �!��U  p"This_stuffs_This_stuffs_ �U  0%��U  �3��U  @'��U   (��U  ���V��  Yst/       Birthday    ����U  ����U  0�Some_stuffs_Some_stuffs_ �U  0���U  ����U  p���U  0���U  ٮnW��  7�t/       Meeting     �g��U  �h��U  pjThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �o��U  �>uW��  �t/       Some_stuffs ���U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  L!"���  !D/      Some_stuffs ����U  ���U  гThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  p���U  �)6���  BI/       Meeting      +��U  �+��U  �/Some_stuffs_Some_stuffs_ �U  �9��U  �:��U  �>��U  �?��U  b����  Dg/      Appointment ����U  `���U   �This_stuffs_This_stuffs_ �U  ����U  `���U  ����U  `���U  �C���  J�/       Some_stuffs ����U  P���U  �Some_stuffs_Some_stuffs_ �U  P���U  ����U  ����U  P���U  �G���  �/      Some_stuffs P��U  ��U  �justforfun_justforfun_ ��U  �"��U  p#��U  p��U  0��U  ��I���  ׏/       Workout ffs ����U  p���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  i�`���  ��/       Meeting ffs �,��U  �-��U  @.This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   3��U  0����  ^�/       Appointment  ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  `���U   ���U  ����U  ��t���  b�/       Workout                        justforfun_justforfun_                                       !����  T�/       Some_stuffs �f��U  �g��U  `hSome_stuffs_Some_stuffs_ �U  `k��U   l��U  �l��U  `m��U  �$����  ��/      Birthday U  P���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  �����  \�/      Birthday                       This_stuffs_This_stuffs_                                     �����  �/       Some_stuffs ����U  P���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  zI/���  �/       Some_stuffs �9��U  �:��U  �>This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  @Q��U  �c����  �-�/       Workout     ����U  ����U  p�Some_stuffs_Some_stuffs_ �U  ����U  @���U  ����U  ����U  �泄��  .�/       Appointment ����U  0���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ���  �1�/       Workout �U  0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  ��ń��  �2�/      Appointment ����U  0���U  ��Some_stuffs_Some_stuffs_ �U  ����U  p���U  0���U  ����U  ,)O���  �U�/      Some_stuffs ���U  ����U  P�justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ����U  �$���  z}�/      Some_stuffs ����U  @���U  ЋSome_stuffs_Some_stuffs_ �U  ����U  `���U   ���U  ����U  HAy���  ��/       Meeting �U   a��U  �a��U  @bSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �f��U  l�z���  q��/       Some_stuffs ���U  ����U  �justforfun_justforfun_ ��U  P���U  ����U  P���U  ���U  )����  ���/       Birthday    �"��U  p#��U  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0��U  �鑆��  m��/       Appointment ���U  0 ��U  � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0&��U  �M����  Ȩ�/      Meeting      ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  P���U  ���U  й��U  �m���  �ƀ/       Appointment ����U  `���U   �Some_stuffs_Some_stuffs_ �U   ���U  ����U  ����U  0��U  �g���  Xʀ/       Appointment  ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  p���U  ���U  ж��U  r���  �ˀ/       Birthday U  ����U  p���U  ��justforfun_justforfun_ ��U  p���U  ����U  ����U  0���U  �����  �ˀ/       Workout �U   ���U  ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �䢇��  O�/      Workout ffs �|��U  �}��U  0~justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  `���U  �ޣ���  ��/       Meeting ffs ����U  ����U  @�This_stuffs_This_stuffs_ �U  ����U   ���U  ����U  `���U  
s����  ��/       Workout     p���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �J����  ���/       Appointment �z��U  `{��U   |Some_stuffs_Some_stuffs_ �U  p��U  0���U  ����U  ����U  �ɼ���  ��/       Appointment ���U  ����U  @�Some_stuffs_Some_stuffs_ �U  `���U  ����U  `���U  ����U  �|O���  ~�/      Workout     P���U  Т��U  ��This_stuffs_This_stuffs_ �U  ���U  ����U  `���U   ���U  4�ֈ��  "=�/      Birthday     E��U  �F��U  0Kjustforfun_justforfun_ ��U  �U��U  �V��U  P[��U  \��U  �����  /A�/       Some_stuffs p?��U  �?��U  p@This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  �D��U  �m���  pC�/       Appointment p;��U  �;��U  P=This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �A��U  ��o���  Ed�/       Appointment ����U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  Z�u���  �e�/       Some_stuffs  ���U  p���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  \q}���  �g�/      Meeting �U   o��U  �o��U  �pSome_stuffs_Some_stuffs_ �U  Ps��U  t��U  �t��U  �u��U  �v~���  h�/       Meeting      %��U  �%��U  @&justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  *��U  ��~���  h�/       Meeting     0��U  ���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0 ��U  3�����  �h�/       Some_stuffs �/��U  p0��U  �4This_stuffs_This_stuffs_ �U  �>��U  �?��U   E��U  �F��U  T}���  v��/      Appointment                    This_stuffs_This_stuffs_                                     r�����  流/       Workout ffs  ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  �����  ���/       Appointment ��U  ���U  �This_stuffs_This_stuffs_ �U  ���U  ���U  p��U  0��U  흿���  E��/      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             $k<���  8ځ/      Appointment ����U  p���U  0�justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  ����U  !HT���  T��/       Appointment �6��U   7��U  �7justforfun_justforfun_ _ �U  P9��U  �9��U  p:��U  0;��U  h�ы��  q �/       Birthday U  0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  ��k���  �'�/      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �{���  �+�/       Some_stuffs ����U  p���U  0�Some_stuffs_Some_stuffs_ �U  ����U  0���U  ���U  ����U  �C���  �O�/       Workout ent 05��U  �5��U  06This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  �:��U  �#���  �Q�/      Some_stuffs ����U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  �m����  nx�/       Appointment �7	��U   8	��U  �8	This_stuffs_This_stuffs_ �U  �:	��U  `;	��U  <	��U  �<	��U  �����  �x�/      Workout     ���U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  1�׎��  �Ƃ/       Appointment pz��U  0{��U  �{Some_stuffs_Some_stuffs_ �U  0~��U  ����U  `���U  ����U  |����  ʂ/      Birthday U  0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  BXp���  ��/       Workout     ����U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  yly���  ��/       Appointment  ��U  ���U  `oSome_stuffs_Some_stuffs_ �U  0r��U  �r��U  �s��U  pt��U  ,~���  -�/      Appointment p��U  0��U  0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p0��U  �c����  �/       Some_stuffs ����U  p���U  ��Some_stuffs_Some_stuffs_ �U  p���U  ����U  ����U  p���U  �����  ��/       Appointment �H��U  pI��U  �IThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �M��U  �����  G�/      Appointment A	��U  �A	��U  PB	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  PF	��U  J�����  �=�/       Some_stuffs ���U  ����U  0�justforfun_justforfun_ ��U  ����U  0���U  ����U  0���U  �w����  �>�/       Some_stuffs p:��U  0;��U  �;Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �?��U  ������  �>�/       Workout     ���U  ����U  P�This_stuffs_This_stuffs_ �U  ���U  ����U  ����U  P���U  j�+���  1_�/       Some_stuffs �m��U  @n��U   oSome_stuffs_Some_stuffs_ �U  �w��U  �x��U  Ps��U  t��U  �<=���  �c�/       Some_stuffs 0f��U  �g��U  �iSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �t��U  �XF���  �e�/      Meeting     P���U  ���U  лThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  ځϑ��  ��/       Workout     ���U  ����U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0���U  ��Ց��  ���/       Meeting      ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  Sߑ��  ��/       Birthday U  @&��U  �&��U  @'justforfun_justforfun_ ��U  p)��U  *��U  �*��U  P+��U  T���  *��/       Birthday    0=��U  �=��U  0>Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �A��U  �����  ���/      Birthday     ���U  ����U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  ��{���  +��/       Workout     ����U  `���U  ��This_stuffs_This_stuffs_ �U   ���U  ����U   ���U  ����U  |3���  _؃/      Meeting     0���U  ����U  p�Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   ���U  �����  ?��/       Workout     е��U  ����U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �ɰ���  F��/      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             (F���  ���/      Appointment е��U  ����U  �Some_stuffs_Some_stuffs_ �U  ����U  ����U  ���U  ����U  ��^���  į�/       Appointment @��U   ��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �i���  ���/       Meeting     Ps��U  t��U  �tThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   z��U  Ox޽��  �Ў/      Meeting     ����U  p���U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0���U  l����  Qю/       Birthday                       Some_stuffs_Some_stuffs_                                     �2���  :Ҏ/       Appointment ����U  ����U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  i����  ֎/       Workout     ����U   ���U  ��This_stuffs_This_stuffs_ �U  @��U   ��U  ���U  @��U  ����  �֎/       Appointment `���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  ���U  Т��U  P���U  ������  �׎/       Meeting     ���U  ����U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  h����  q��/       Some_stuffs 0���U  ����U  p�justforfun_justforfun_ ��U  P
��U  �
��U  @���U  ����U  �����  ��/       Meeting ffs 0���U  ����U  0�This_stuffs_This_stuffs_ �U  ����U  0���U  ���U  ����U  �����  �!�/      Some_stuffs ���U  ����U  0�justforfun_justforfun_ ��U   ���U  ����U  ����U  @���U  ��#���  �#�/       Workout     ���U  ����U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  I�����  �H�/       Appointment P��U  ���U  PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p#��U  ������  oJ�/       Birthday    ����U  P���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  -˿��  �N�/      Some_stuffs � ��U  �!��U  p"Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   (��U  �aE���  �m�/       Workout ent �z��U  P{��U  |This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  �J���  ?o�/       Some_stuffs 0f��U  �g��U  �iSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �t��U  �*X���  �r�/      Appointment ���U  ����U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  @�]���  (t�/       Birthday    p���U  0���U  ��Some_stuffs_Some_stuffs_ �U  ����U  ����U   ���U  ����U  ������  ���/       Birthday                       justforfun_justforfun_ _                                     �L����  ���/      Meeting     ���U  ����U  P�This_stuffs_This_stuffs_ �U  г��U  p���U  p���U  0���U  ᱅���  쿏/       Meeting ent `���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  `���U  ����U  ����U  �ʈ���  ���/       Meeting     ��U  ���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0��U  �����  z�/       Meeting     06��U  �6��U  p7justforfun_justforfun_ ��U  �9��U  �:��U  p;��U  �;��U  �����  ]�/      Workout     ����U  @���U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  �P����  ��/       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             LM����  �W�/      Appointment ����U  ����U   �This_stuffs_This_stuffs_ �U  Ћ��U  ����U   ���U  ����U  �����  �X�/       Birthday    ����U  p���U  0�This_stuffs_This_stuffs_ �U  ���U  ����U  ����U  @���U  �����  AZ�/       Meeting     ����U   ���U  ��justforfun_justforfun_ _ �U  ����U  `���U   ���U  ���U  �i����  Æ�/       Workout     `\��U  �\��U  �]Some_stuffs_Some_stuffs_ �U  �_��U  p`��U  �`��U  �a��U  t�����  ʆ�/      Meeting      ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  `���U   ���U  ����U  �B���  ��/       Meeting     �G��U   H��U  �HSome_stuffs_Some_stuffs_ �U  �J��U  @K��U  �K��U  @L��U  �<���  Ъ�/       Workout ent ���U  0��U  �justforfun_justforfun_ ��U  ���U  ���U  p��U  0��U  �����  x��/       Birthday    p��U  0��U  0justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  p0��U  T$���  ��/      Birthday U   ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  Dn����  l͐/      Appointment �>��U  ?��U  �?This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �D��U  �cM���  0��/      Birthday nt �z��U  P{��U  |justforfun_justforfun_ _ �U  �~��U  P��U  ���U  P���U  �h����  ��/      Appointment е��U  ����U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �=����  !�/       Birthday nt  ���U  ����U  `�This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  ����U  
(i���  �A�/       Meeting �U  0���U   ���U  @�This_stuffs_This_stuffs_ �U  p���U  0���U  ����U  `���U  ��u���  	E�/      Meeting     P���U  ����U  P�Some_stuffs_Some_stuffs_ �U  ����U  p���U  ����U  ����U  +i����  �G�/       Some_stuffs 0f��U  �g��U  �iSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �t��U  �x����  �G�/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_              �����  �J�/       Some_stuffs                    Some_stuffs_Some_stuffs_                                     UM���  vp�/      Workout     ���U  ����U  ��justforfun_justforfun_ ��U  ����U  @���U  0���U   ���U  0f ���  �p�/       Some_stuffs `k��U   l��U  �lThis_stuffs_This_stuffs_ �U  `o��U   p��U  �p��U  �q��U  ������  a��/       Workout     p���U  0���U  ��justforfun_justforfun_ ��U  p���U  ����U  ����U  0���U  ͢���   ��/       Birthday    �Q��U   R��U  �RThis_stuffs_This_stuffs_ �U  �T��U  `U��U   V��U  �V��U  ������  3��/      Birthday    ����U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �
��U  �^����  d��/       Appointment                    justforfun_justforfun_                                        I5���  ���/       Birthday    ����U  P���U   �Some_stuffs_Some_stuffs_ �U  ���U  А��U  ����U  p���U  �@���  ���/      Some_stuffs ����U  ����U  `�Some_stuffs_Some_stuffs_ �U   ���U  ���U  ����U  ���U  |�v���  �	�/      Some_stuffs ����U  ����U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  1�����  ~�/       Workout     Ѕ��U  ����U  �justforfun_justforfun_ ��U  ����U  P���U  ���U  Ћ��U  ������  ,�/      Workout     �g��U  �h��U  pjSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �o��U  1�����  T�/       Meeting �U  ����U  `���U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  b]����  V�/       Some_stuffs p���U  0���U  ��This_stuffs_This_stuffs_ �U  p���U  ����U  ����U  0���U  �����  Z�/       Workout     ����U  @���U  ��justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  ���U  +*����  iZ�/       Appointment p���U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  xj����  �Z�/       Appointment е��U  ����U  �Some_stuffs_Some_stuffs_ �U  ����U  ����U  ���U  ����U  ŗ=���  \~�/      Workout �U  0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  ��>���  �~�/       Appointment ����U  ����U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ������  ϥ�/      Some_stuffs ���U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  �7a���  ɒ/       Meeting      ��U  ���U   Some_stuffs_Some_stuffs_ �U  @!��U  �!��U  @"��U   #��U  |�v���  Β/      Appointment ����U  ����U  ��justforfun_justforfun_ ��U  ����U  p���U  0���U  ����U  �Oy���  /ϒ/       Meeting     0���U  ����U  ��justforfun_justforfun_ ��U  p���U  0���U  ����U  ����U  @���  ���/       Meeting     0���U  ����U  ��Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  p���U  ��I���  ŝ/      Appointment p���U  0���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  �f����  ��/       Meeting     ����U  `���U  �Some_stuffs_Some_stuffs_ �U  p���U  ����U  ����U  0���U  �� ���  ��/      Appointment ����U  ����U  p�This_stuffs_This_stuffs_ �U  ����U  @���U  ����U  ����U  ����  :��/       Some_stuffs ���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �&y���  ��/       Appointment `���U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  E�}���  ��/      Some_stuffs ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Т��U  �����  ��/       Meeting     PH��U  I��U  �Ijustforfun_justforfun_ ��U  PL��U  M��U  �M��U  �N��U  %<����  �`�/       Workout     �~��U  P��U  �This_stuffs_This_stuffs_ �U  ���U  ����U  ���U  Ѓ��U  t^����  fb�/       Workout     ����U  P���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ������  �d�/       Some_stuffs л��U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  �\����  �e�/      Meeting      ��U  ���U  @ This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �$��U  *]����  Ih�/       Appointment ���U  ���U  pThis_stuffs_This_stuffs_ �U   &��U  �&��U  0��U  ���U  ������  dh�/       Appointment �i��U  pj��U  0kThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  po��U  �tF���  ҈�/      Workout                        justforfun_justforfun_                                       ��I���  ���/       Birthday    �y��U   z��U  �zSome_stuffs_Some_stuffs_ �U  �}��U  `~��U   ��U  ���U  �`���  b��/       Birthday    @���U  ���U  p�Some_stuffs_Some_stuffs_ �U  д��U  P���U  ���U  ж��U  ������  g��/      Workout     ���U  ����U  0�justforfun_justforfun_ ��U   ���U  ����U  ����U  @���U  @����  �۞/       Some_stuffs pG��U  �G��U  �HSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pL��U  �����  /��/       Birthday    �$	��U  `%	��U  &	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   *	��U  \����  ���/      Some_stuffs ����U  ����U  p�This_stuffs_This_stuffs_ �U  0���U  ����U  0���U  ����U  Qv���  ��/       Birthday    ����U  ���U  ��This_stuffs_This_stuffs_ �U  ����U  ���U  ����U  ���U  �����  w(�/       Appointment @X��U  �X��U  �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ^��U  p�����  �)�/       Birthday U  `V��U   W��U  �WThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U   ]��U  F�����  l*�/      Some_stuffs p���U  0���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  �8����  �u�/      Some_stuffs p���U  0���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  Y����  �z�/       Some_stuffs ����U  ����U  p�justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ����U  �}���  �/      Meeting      b��U  �b��U   cSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �g��U  0z  �  >ş/       Meeting ent P���U  ����U  P�Some_stuffs_Some_stuffs_ �U  ����U  P���U  ����U  P���U  �++  �  �ɟ/       Workout     ���U  ���U  pThis_stuffs_This_stuffs_ �U   &��U  �&��U  0��U  ���U  uO�  �  
�/      Appointment  ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  `���U   ���U  ����U  ��  �  *�/       Meeting                        This_stuffs_This_stuffs_                                     �e: �  ��/      Some_stuffs 0f��U  �g��U  �iThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �t��U  ��L �  ��/       Some_stuffs @���U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @	��U  y�L �  ��/       Workout �U  ���U  ����U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  r<� �  &9�/       Some_stuffs �	��U  @	��U  �	Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  @	��U  p�� �  f<�/       Meeting �U  ����U  p���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  ��� �  �=�/      Birthday    @.��U  �.��U  �/Some_stuffs_Some_stuffs_ �U  �2��U   3��U   4��U  �4��U  ��z �  a�/      Workout      ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��| �  ya�/       Some_stuffs  ��U  ���U  @Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ,& �  ͌�/      Workout     ����U  @���U  �This_stuffs_This_stuffs_ �U  P���U  ���U   ���U  ����U  �)� �  ��/       Meeting     �`��U  `a��U   bThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `f��U  �J� �  歠/      Some_stuffs @p��U   q��U   �Some_stuffs_Some_stuffs_ �U  @t��U  �t��U  �u��U  v��U  XN� �  筠/       Workout     ���U  ж��U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  }� �  ʱ�/       Some_stuffs p��U  0��U   &Some_stuffs_Some_stuffs_ �U  ���U  p��U  0��U  ���U  HQ �  ]٠/       Appointment @��U  ���U  @justforfun_justforfun_ _ �U  @��U  ���U  @��U   ��U  0�� �  ���/       Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             Eq� �  L��/      Some_stuffs �Q��U  PR��U  �RSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  `r��U  �Sh �  � �/       Appointment PF��U  �F��U  PGjustforfun_justforfun_ ��U  �I��U  �J��U  K��U  �K��U  *� �  �&�/       Appointment ����U   ���U  ��justforfun_justforfun_ ��U  @���U  ����U  @���U  ����U  �^� �  )�/       Birthday    ���U  p���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �] �  K�/      Workout �U  ��	��U   �	��U  Ё	Some_stuffs_Some_stuffs_ �U  0�	��U  ��	��U  0�	��U  ��	��U  ��� �  8n�/       Workout     ���U  ����U  �justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ���U  \<� �  �n�/       Meeting     P���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  P���U  ���U  ����U  3� �  �p�/       Workout     �I��U  �J��U  KThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �O��U  � �  .r�/      Birthday    p���U  ����U  p�Some_stuffs_Some_stuffs_ �U  0���U  ����U  p���U  ����U  j	� �  qr�/       Meeting     �}��U  ~��U  �~This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  �LG �  x��/       Some_stuffs p��U  0��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p��U  ��� �  ���/       Workout     @���U  ����U  @�Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  �� �  ���/      Meeting      ��U  ���U   justforfun_justforfun_ ��U  @��U  ���U  @��U  ���U  �� �  L��/       Meeting     �|��U  p}��U  �}This_stuffs_This_stuffs_ �U  ���U  ����U  ���U  Ё��U  ��	 �  ��/       Some_stuffs p ��U  0��U  pSome_stuffs_Some_stuffs_ �U  0��U  ���U  p��U  0��U  �2	 �  ��/      Some_stuffs  ���U  ���U  ��Some_stuffs_Some_stuffs_ �U  ���U  ����U  P���U  ���U  !��	 �  �7�/       Workout     @���U  ����U  @�This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  @���U  <�	 �  79�/      Birthday    ����U  p���U  �This_stuffs_This_stuffs_ �U  ����U  0���U  ����U  p���U  �r0
 �  :Z�/      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �1
 �  �Z�/       Workout     �P��U  Q��U  �Qjustforfun_justforfun_ ��U  T��U  �T��U  PU��U  �U��U  ���3 �  �	�/      Some_stuffs P��U  ���U  PThis_stuffs_This_stuffs_ �U  ���U  �	��U  �"��U  p#��U  (��3 �  	�/       Workout     ���U  p��U  0This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  �}4 �  ^.�/      Birthday    `���U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  )=�4 �  I4�/       Appointment p��U  ���U  �justforfun_justforfun_ ��U  p��U  0��U  ���U  p��U  ���5 �  ��/       Appointment  ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  `���U  ����U  `���U  ���5 �  ���/      Some_stuffs  ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  }H6 �  ߣ�/      Appointment 0���U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0���U  B�_6 �  詭/       Some_stuffs P���U  ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  ��b6 �  ���/       Appointment @^��U  �^��U  �OSome_stuffs_Some_stuffs_ �U  pR��U  �R��U  �S��U  pT��U  ��6 �  �ѭ/      Birthday    0���U  ����U  p�justforfun_justforfun_ ��U  ����U   ���U  @���U   ���U  <��7 �  w��/      Workout     p��U  0��U  0Some_stuffs_Some_stuffs_ �U   +��U  �+��U  �/��U  p0��U  "&�7 �  ��/       Birthday    P���U  ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  A��7 �  ���/       Appointment �9��U  �:��U  p;justforfun_justforfun_ ��U  �>��U  ?��U  �?��U  P@��U  O�8 �  A�/      Birthday    ����U  ���U  ��Some_stuffs_Some_stuffs_ �U  ����U  ���U  ����U  ���U  ʌ8 �  M�/       Some_stuffs ����U  `���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  o!8 �  
�/       Some_stuffs ����U  `���U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0��U  8�!8 �  �/       Some_stuffs ����U  p���U  0�Some_stuffs_Some_stuffs_ �U  ����U  ����U  p ��U  0��U  ��!8 �  %�/       Birthday    �w��U  �x��U  PsSome_stuffs_Some_stuffs_ �U  v��U  �v��U  0~��U  �~��U   ��8 �  @E�/       Some_stuffs @���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  )��8 �  �F�/       Birthday    �d��U  �e��U  @fThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @j��U  ��D9 �  �g�/       Some_stuffs ����U  ����U  НSome_stuffs_Some_stuffs_ �U  0���U  ���U  p���U  0���U  �c9 �  ]o�/      Birthday    �f��U  �g��U  `hSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `m��U  �=�9 �  I��/      Meeting                        Some_stuffs_Some_stuffs_                                     �~: �  ѷ�/      Birthday nt ����U  ���U  ��justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  @���U  ɤ�: �  M��/       Workout  U  ����U  P���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  Z�: �  缮/       Meeting ffs �w	��U  `x	��U  �x	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �|	��U  ��; �  �߮/      Birthday                       Some_stuffs_Some_stuffs_                                     �E; �  �/       Some_stuffs @'��U  �'��U  @(justforfun_justforfun_ ��U  �*��U  P+��U  �+��U  �,��U  �"; �   �/       Appointment �*��U  p+��U  0,justforfun_justforfun_ ��U  �.��U  p/��U  00��U  �0��U  4��; �  ��/      Meeting �U  �,��U  �-��U  @.Some_stuffs_Some_stuffs_ �U   1��U  �1��U  �2��U   3��U   9J< �  �-�/       Meeting     ���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �O< �  �.�/      Workout     ����U  `���U  ��justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ���U  ���< �  /U�/       Some_stuffs �w��U  px��U  0yjustforfun_justforfun_ ��U  �{��U  0|��U  �|��U  �}��U  �t�< �  �V�/      Some_stuffs Ѕ��U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Ћ��U  @��= �  h��/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ���= �  /      Workout     ����U  0���U  P
Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  ��$> �  ��/       Meeting  nt �X��U  @Y��U  �YThis_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  @^��U  �0(> �  ���/      Birthday    ���U  p��U  0This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  !�9? �  ��/       Appointment Р��U  ����U  P�justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ����U  �CQ? �  	��/      Workout     ���U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ���? �  :�/      Birthday fs 0��U  ���U  0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �<��U  ��? �  ��/       Birthday    @\��U   ]��U  �]This_stuffs_This_stuffs_ �U  �`��U  `a��U   b��U  �b��U  ��z@ �  7@�/       Workout     x��U  �x��U  �yjustforfun_justforfun_ ��U  |��U  �|��U  �}��U  ~��U  J~@ �  A�/      Appointment ����U  @���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  	�A �  �f�/       Birthday    ���U  ����U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �A �  j�/       Some_stuffs `���U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `���U  hX�A �  щ�/       Appointment �z��U  `{��U   |Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  A�A �  ��/       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �q�A �  D��/       Meeting     �<��U  �=��U   >This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �A��U  x>B �  ճ�/       Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             sEB �  ���/       Some_stuffs  $��U  �%��U   +justforfun_justforfun_ ��U  �4��U  p5��U  �9��U  �:��U  R*IB �  ���/       Some_stuffs  ���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  U�LB �  v��/      Birthday    ����U  `���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  H`�B �  }۰/       Some_stuffs �.��U  p/��U  00Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �4��U  �^�B �  �ް/      Birthday    0���U  ����U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  [�bC �  ���/       Appointment ��U  ���U  Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  P��U  �eC �  `��/       Appointment ����U  ����U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��tC �  K�/       Appointment ����U  p���U  0�This_stuffs_This_stuffs_ �U  ���U  ����U  ����U  @���U  ���C �  �/      Some_stuffs p7��U  08��U  �8Some_stuffs_Some_stuffs_ �U  p;��U  �;��U  P=��U  >��U  ͂D �  (�/      Meeting     P���U  ����U  @This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  H�D �  )�/       Birthday    p��U  0��U  �Some_stuffs_Some_stuffs_ �U  ���U  ���U  p��U  ���U  ,#5E �  v�/      Some_stuffs ����U  @���U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  QGGE �  �z�/       Meeting �U  ����U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  ��o �  �K�/       Workout      ��U  ���U   This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  �/�o �  �P�/       Meeting     ���U  ����U  P�justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  P���U  �J�o �  �Q�/      Meeting ent @g��U  �g��U  �hThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   m��U  `^p �  �p�/       Some_stuffs `���U   ���U  ��Some_stuffs_Some_stuffs_ �U  `���U   ���U  ����U  `���U  #�p �  Tq�/       Birthday     ���U  ����U  `�Some_stuffs_Some_stuffs_ �U  ����U  `���U  `���U   ���U  �*p �  lu�/       Workout �U  �v��U  �w��U  xSome_stuffs_Some_stuffs_ �U  �z��U  P{��U  |��U  �|��U  ͋3p �  �w�/      Workout     �p��U  �q��U  0rSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0w��U  :ȼp �  Ӛ�/       Some_stuffs ����U  p���U  0�This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  @���U  )��p �  	��/       Some_stuffs  Z	��U  �Z	��U   [	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �^	��U  (��p �  )��/       Appointment ����U  `���U   �Some_stuffs_Some_stuffs_ �U  ����U  ���U  ����U  ���U  5Oq �  b��/      Birthday    Ю��U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  ��Oq �  d��/       Birthday    p��U  0��U  �This_stuffs_This_stuffs_ �U  ���U  ���U  p��U  ���U  �~�q �  �/       Workout      ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  ���q �  ��/       Appointment ����U  ����U   �justforfun_justforfun_ ��U  Н��U  p���U  0���U  ����U  ���q �  �/       Workout     ����U  @���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �I�q �  �/      Meeting     ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  @���U  0���U   ���U  ��r �  $�/       Appointment  ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  D+�r �  ��/      Some_stuffs  ���U  ����U  ��This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ж��U  R�#s �  28�/       Some_stuffs P	��U  �	��U  �	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0!	��U  ��)s �  �9�/       Birthday    ����U  ����U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��/s �  S;�/      Appointment                    This_stuffs_This_stuffs_                                     �o�s �  X_�/       Birthday    ����U  p���U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  ���s �  �_�/       Meeting      :��U  �:��U  0;This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �>��U  ��_t �  1��/      Birthday    @'��U   (��U  �(justforfun_justforfun_ ��U  �+��U   ,��U  �,��U  �-��U   ��t �   ��/       Meeting     ����U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  q��t �  &��/       Some_stuffs pA��U  �A��U  pBThis_stuffs_This_stuffs_ �U  �D��U  @{��U  0F��U  �F��U  �t �  `��/       Birthday    @_��U  P���U  �`justforfun_justforfun_ ��U  �b��U  @c��U  �c��U  �d��U  ���t �  G��/      Appointment  b��U  �b��U   cjustforfun_justforfun_ _This_stuffs_This_stuffs_ �U  �g��U  ��vu �  �н/       Meeting ffs ����U  p���U  0�This_stuffs_This_stuffs_ �U  0���U  ���U  p���U  ���U  h߄u �  1Խ/       Workout     ����U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ]t�u �  �׽/      Some_stuffs ����U  p���U  �justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  ���U  ZRv �  g��/       Workout ffs P���U  ����U  P�justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  P���U  �cv �  0��/       Some_stuffs  ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��v �  ���/      Some_stuffs ���U  ����U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  ��v �  ���/       Workout ffs ����U  p���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  ��v �  ��/       Appointment ����U  `���U   �This_stuffs_This_stuffs_ �U   ���U  ����U  ����U   ���U  R��v �  � �/       Meeting     P���U  ����U  ��justforfun_justforfun_ _ his_stuffs_This_stuffs_ �U  P���U  ���v �  �"�/      Appointment T��U  �T��U  PUjustforfun_justforfun_ ��U   W��U  �W��U  @X��U  �X��U  �v �  U#�/       Appointment л��U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  ��Ow �  �I�/      Birthday U  `���U   ���U  ��justforfun_justforfun_ ��U  `���U   ���U  ����U  `���U  �Sw �  �J�/       Birthday    ���U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  ص�w �  �q�/       Appointment ���U  ���U  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0��U  ��zx �  +��/       Some_stuffs �[��U  `\��U  �\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @a��U  �
�x �  䚾/       Meeting ent ����U  @���U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  bh
y �  ���/       Appointment �C��U  �D��U  EThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  I��U  i�y �  ���/       Meeting ffs ���U  ���U  pSome_stuffs_Some_stuffs_ �U  p��U  0��U  ���U  ���U  ;�y �  ���/       Some_stuffs  !��U  �!��U  `"Some_stuffs_Some_stuffs_ �U  �$��U   %��U  �%��U   &��U  ��y �  ���/       Some_stuffs P[��U  \��U  �`This_stuffs_This_stuffs_ �U   l��U  �l��U  �g��U  �h��U  щ�y �  B�/       Appointment `���U   ���U  НSome_stuffs_Some_stuffs_ �U  0���U  ���U  ����U  p���U  l��y �  �/      Workout     �P��U  @Q��U  �UThis_stuffs_This_stuffs_ �U  �`��U  �a��U  `f��U   g��U  Y7=z �  �	�/       Birthday    |��U  �|��U  �}justforfun_justforfun_ ��U  ���U  P���U  ���U  ����U  ��Dz �  z�/      Workout                        justforfun_justforfun_                                       3Qz �  ��/       Appointment �`��U  �a��U  `fThis_stuffs_This_stuffs_ �U  �g��U  �h��U  pj��U  0k��U  �Vz �  
�/       Workout     `���U  ���U  ��Some_stuffs_Some_stuffs_ �U  ����U  ���U  ����U  ���U  �Xz �  ��/       Appointment @*��U   +��U  �+Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @0��U  ��Yz �  ��/       Meeting     ���U  ���U  0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @��U  ��z �  A/�/       Some_stuffs  9��U  �9��U  `:Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �>��U  Z�z �  G5�/       Appointment p���U  ����U  ��justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  p���U  ��z �  D7�/      Some_stuffs ����U  P���U  �Some_stuffs_Some_stuffs_ �U  `���U   ���U  ���U  ����U  �m{ �  OW�/       Birthday    �B��U  pC��U  �CThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   H��U  ��q{ �  xX�/       Birthday U  ����U  @���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��~{ �  �[�/       Birthday    ����U  p���U  0�This_stuffs_This_stuffs_ �U  0���U  ����U  p���U  0���U  �^| �  邿/      Workout     �)��U  0*��U  �*justforfun_justforfun_ ��U  p-��U  0.��U  �.��U  p/��U  ):| �  i��/       Appointment �T	��U  @U	��U  �U	This_stuffs_This_stuffs_ �U  �W	��U  @X	��U  �X	��U  pY	��U  �N�| �  ���/       Meeting     �_��U  �`��U   ajustforfun_justforfun_ _ �U  �c��U  @d��U  �d��U  �e��U   @} �  �ο/      Appointment �y��U  Pz��U  �zThis_stuffs_This_stuffs_ �U  �}��U  ~��U  �~��U  P��U  0fG} �  �п/       Appointment p���U  ����U  ��Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ����U  ��} �  ���/      Workout     P���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  P���U  ���U  ����U  Ćd~ �  ��/      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_              � �  �C�/       Meeting �U  P[��U  \��U  �`Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �h��U  �r �  �D�/       Some_stuffs �G��U  0H��U  �HThis_stuffs_This_stuffs_ �U  �K��U  0L��U  �L��U  �M��U  Y� �  �H�/       Appointment P[��U  \��U  �`This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �h��U  6$ �  �I�/      Meeting      2��U  �2��U   3This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   7��U  q�� �  �j�/       Workout     PO��U  �O��U  �PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �T��U  <�� �  7l�/      Appointment @���U  ����U  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �L� �  vp�/       Birthday    ����U  ����U  НSome_stuffs_Some_stuffs_ �U  0���U  ���U  p���U  0���U  h�K� �  q��/       Workout     ���U  ����U  p�justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  P���U  �y΀ �  ��/       Birthday    `_��U   `��U  �`Some_stuffs_Some_stuffs_ �U   c��U  �c��U  `d��U  �d��U  L�Ԁ �  ���/      Meeting     ����U  p���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  �*b� �  ���/      Workout     P���U  ����U  @This_stuffs_This_stuffs_ �U  ����U  ����U  p���U  ����U  y�e� �  ���/       Birthday    �W��U  �X��U  @YThis_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  �n��U  ��[(�  �T
 /      Birthday    ����U  @���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  i8_(�  �U
 /       Appointment  ��U  ���U  �This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  �%��U  ���(�  :y
 /      Workout     ����U  ����U  Нjustforfun_justforfun_ ��U  0���U  ���U  p���U  0���U  [��(�  '}
 /       Appointment �/��U  @0��U   1Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �5��U  hl�(�  Q~
 /       Workout     �g��U  �h��U  pjSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �o��U  �� )�  8
 /       Meeting      ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  `���U  ����U  `���U  �[�)�  ֟
 /       Birthday fs  ��U  ���U   This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ��U  ㍆)�  l�
 /       Some_stuffs �1��U   2��U  �2Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P7��U  �<�)�  "�
 /       Some_stuffs @*��U   +��U  �+This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  @0��U  �D�)�  ��
 /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �*�  ��
 /       Some_stuffs ����U  ����U  `�This_stuffs_This_stuffs_ �U  ����U  0���U  ����U  P���U  ��%*�  <�
 /      Some_stuffs ���U  ����U  ��justforfun_justforfun_ ��U  ����U  @���U  0���U   ���U  �e4*�  ��
 /       Appointment ����U  ����U  p�This_stuffs_This_stuffs_ �U  ����U  @���U  ����U  ����U  ]R�*�  k�
 /      Some_stuffs ����U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  Hz�*�  ��
 /       Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             Jٽ*�  �
 /       Appointment ����U  `���U  ��This_stuffs_This_stuffs_ �U  ����U  `���U  е��U  ����U  z#W+�  [ /       Appointment ����U  � ��U  @Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  �#W+�  [ /      Birthday    ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  F[+�  j /       Workout �U  @��U  ���U  @Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   ��U  c+�  j /       Meeting �U  и��U  ����U  P�Some_stuffs_Some_stuffs_ �U  м��U  P���U  ���U  о��U  �k+�  � /       Appointment е��U  ����U  �This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  ����U  ���+�  �B /       Appointment ����U  `���U  ��justforfun_justforfun_ ��U   ���U  ����U  `���U  ����U  a~,�  �D /       Meeting     �>��U  ?��U  �?This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �D��U  ��{,�  Oc /      Meeting     ���U  ����U  0�Some_stuffs_Some_stuffs_ �U   ���U  ����U  ����U  @���U  �Y-�  � /       Some_stuffs  ��U  ���U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  �-�  �� /       Workout      ��U  ���U  0justforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U  ���U  mu"-�  � /       Workout     P	��U  �	��U  �	justforfun_justforfun_ _ �U  �	��U  @	��U  �	��U  @	��U  �+-�  $� /       Some_stuffs  E��U  �F��U  0KThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  \��U  
O+-�  5� /       Birthday    ����U  0���U  ��Some_stuffs_Some_stuffs_ �U  ����U  p���U  0���U  ����U  ��0-�  �� /      Workout      o��U  �o��U  �pjustforfun_justforfun_ ��U  Ps��U  t��U  �t��U  �u��U  Ľ�-�  � /      Some_stuffs �m��U  @n��U   oSome_stuffs_Some_stuffs_ �U  �w��U  �x��U  Ps��U  t��U  (6K.�  �� /       Some_stuffs  E��U  �F��U  0KSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  \��U  'X.�  9� /      Some_stuffs �2��U   3��U   4Some_stuffs_Some_stuffs_ �U  `6��U   7��U  �7��U  `8��U  L0Y.�  }� /       Appointment  c��U  �c��U  `dThis_stuffs_This_stuffs_ �U  �f��U  �g��U  `h��U   i��U  }�Y.�  �� /       Appointment ���U  ����U  ��justforfun_justforfun_ ��U  ����U  ����U  P���U  ����U  Z.�  �� /       Workout     ����U  @���U  �This_stuffs_This_stuffs_ �U  P���U  ���U   ���U  ����U  Qp\.�  R� /       Meeting �U  ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  @���U  0���U   ���U  q/�.�  � /       Some_stuffs  ���U  ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  ���.�  ) /      Appointment ����U  @���U  P�Some_stuffs_Some_stuffs_ �U  P���U  Т��U  ����U  P���U  \ʁ/�  k) /      Meeting �U  0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  ��0�  �M /      Meeting     ���U  p��U  0Some_stuffs_Some_stuffs_ �U  ���U  0 ��U  � ��U  �!��U  �9'0�  �S /       Appointment �t��U  �u��U  vSome_stuffs_Some_stuffs_ �U  `y��U   z��U  �z��U  `{��U  �s�0�  Wt /       Appointment PI	��U  �I	��U  PJ	justforfun_justforfun_ 	��U  PL	��U  M	��U  �M	��U  N	��U  �g�0�  �u /      Workout      ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  `���U   ���U  ����U  ��0�  w /       Workout     ����U  ���U  ЮThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  ��O1�  �� /       Appointment P���U  ����U  P�justforfun_justforfun_ ��U  ����U  P���U  ���U  ����U  ��`1�  � /       Appointment ���U  ����U  P�This_stuffs_This_stuffs_ �U  ���U  ����U  ����U  P���U  \��1�  �� /      Birthday     ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `���U  ��2�  9� /      Meeting ent ����U  `���U  ��justforfun_justforfun_ _ �U  ���U  `��U  ��U  ���U  ���2�  �� /       Workout     ����U  `���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  1_3�  ^ /       Some_stuffs  ��U  ���U  `oSome_stuffs_Some_stuffs_ �U  0r��U  �r��U  �s��U  pt��U  �*3�   /      Workout     �/��U  p0��U  �4This_stuffs_This_stuffs_ �U  �>��U  �?��U   E��U  �F��U  �Ҩ3�  �9 /       Birthday    ����U  @���U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  I�3�  �9 /       Some_stuffs ���U  p���U  �Some_stuffs_Some_stuffs_ �U  0���U  ���U  p���U  ���U  �ҷ3�  e= /       Birthday    0���U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  {�3�  �> /       Some_stuffs  ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  �jS4�  :e /       Meeting      +��U  �+��U  �/justforfun_justforfun_ ��U  �9��U  �:��U  �>��U  �?��U  ,O�4�  �� /      Some_stuffs `?��U   @��U  �NThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �D��U  9q�4�  s� /       Meeting     00��U  �0��U  p1Some_stuffs_Some_stuffs_ �U  04��U  �4��U  05��U  �5��U  +�x5�  I� /       Workout     ����U  P���U  �Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ����U  �	5�  � /       Workout �U  ����U  ����U  ��justforfun_justforfun_ ��U  ����U  p���U  0���U  ����U  Ъ�5�  � /       Meeting �U  ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  @���U  0���U   ���U  ~��5�  � /      Appointment ���U  ����U  P�Some_stuffs_Some_stuffs_ �U  @���U  ���U  ���U  ����U  c�6�  |� /       Appointment ����U  @���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  �w6�  �� /       Workout     p��U  0��U  �Some_stuffs_Some_stuffs_ �U  ���U  ���U  p��U  ���U  ��6�  �� /       Appointment 0f��U  �g��U  �iSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �t��U  �6�  �� /       Birthday    0���U  ���U  p�justforfun_justforfun_ ��U  ����U  @���U  P���U  ���U  f�!6�  �� /      Workout �U  ����U  0���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  RA�6�  �� /       Appointment ����U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  lG�6�  5� /      Some_stuffs                    This_stuffs_This_stuffs_                                     Q@�6�  R  /       Workout     ����U  P���U  �This_stuffs_This_stuffs_ �U  ����U  `���U  Э��U  P���U  0�W7�  �* /       Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ���7�  �J /       Some_stuffs  ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  `���U  ����U  `���U  r��7�  FM /       Workout     ���U  0��U  �Some_stuffs_Some_stuffs_ �U  p��U  0��U  ���U  0��U  �]�7�  �N /      Some_stuffs 0%��U  �3��U  @'This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ,��U  ���7�  R /       Workout     P[��U  \��U  �`Some_stuffs_Some_stuffs_ �U   l��U  �l��U  �g��U  �h��U  8Gf8�  3p /       Appointment P[��U  \��U  �`justforfun_justforfun_ ��U   l��U  �l��U  �g��U  �h��U  �Yp8�  �r /      Meeting     ����U  ���U  ��This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  P���U  j��8�  �x /       Meeting ent ����U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��9�  Ě /       Meeting ffs p���U  0���U  ��justforfun_justforfun_ ��U  0���U  ����U  p���U  ���U  I�9�  �� /       Workout     0���U  ����U  0�justforfun_justforfun_ ��U  0���U  ���U  ����U  0���U  �O9�  � /       Appointment x��U  �x��U  �ySome_stuffs_Some_stuffs_ �U   |��U  �|��U  �}��U  `~��U  ��9�  ^� /      Meeting     ����U  `���U   �This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U   �9�  4� /       Meeting     ���U  ����U  �Some_stuffs_Some_stuffs_ �U  Ѕ��U  ����U  ���U  ����U  T<:�  v� /      Some_stuffs ����U  P���U  ЪThis_stuffs_This_stuffs_ �U  ����U  ���U  Ю��U  ����U  ��c�  A� /       Some_stuffs ���U  P��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p��U  4u�c�  "� /      Appointment �.��U  p/��U  00justforfun_justforfun_ ��U  �2��U  p3��U  04��U  �4��U  \7�d�  �� /      Workout �U  ����U  P���U  �justforfun_justforfun_ ��U  `���U   ���U  ���U  ����U  ��e�  �� /       Some_stuffs  1��U  �1��U  �2Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   7��U  e�e�  @� /      Appointment 0���U  ����U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��;e�  p� /       Workout     P���U  Щ��U  P�Some_stuffs_Some_stuffs_ �U  p���U  ���U  p���U  0���U  �=e�  �� /       Some_stuffs `_��U   `��U  �`This_stuffs_This_stuffs_ �U   c��U  �c��U  `d��U  �d��U  �)�e�  s /      Appointment ����U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��lf�  }8 /      Birthday U  0f��U  �g��U  �iThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �t��U  :�f�  W /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ���f�  e\ /       Appointment ���U  ���U  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ܇g�  �~ /      Appointment ����U  @���U  �Some_stuffs_Some_stuffs_ �U  P���U  ���U   ���U  ����U  �w�g�  �� /       Some_stuffs ����U  ����U  p�This_stuffs_This_stuffs_ �U  0���U  ����U  0���U  ����U  ���g�  �� /       Some_stuffs 0���U  ����U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0���U  {�g�  [� /       Appointment @f��U  �f��U  @gThis_stuffs_This_stuffs_ �U  �i��U  @j��U   k��U  �k��U  A�h�  ȥ /       Birthday U  �t��U  �u��U  vThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `{��U  �@h�  �� /      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �.,h�  � /       Appointment ����U  P���U  �This_stuffs_This_stuffs_ �U  P���U  ����U  ����U  P���U  �^�h�  �� /       Meeting     p���U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��h�  � /       Birthday     ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  cv�h�  �� /       Meeting �U  (	��U  �(	��U  @)	justforfun_justforfun_ 	��U  �+	��U   ,	��U  �,	��U   -	��U  �C�h�  2� /      Meeting     ����U  0���U  �Some_stuffs_Some_stuffs_ �U  p���U  0���U  ����U  0���U  �Ui�  � /       Meeting     �2��U  p3��U  04justforfun_justforfun_ ��U  06��U  �6��U  p7��U  08��U  3�Vi�  ~� /       Workout ffs �N��U  PO��U  0ASome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �E��U  �ei�  %� /       Some_stuffs ���U  ����U  P�Some_stuffs_Some_stuffs_ �U  @���U  ���U  ���U  ����U  <Ifi�  w� /      Appointment 0���U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  L�gi�  �� /       Workout �U  0f��U  �g��U  �iThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �t��U  ���i�  g /      Workout ffs Р��U  ����U  P�Some_stuffs_Some_stuffs_ �U  ���U  ����U  ���U  ����U  �K�i�  � /       Workout ent ����U  0���U  ��Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ����U  @��i�  � /       Some_stuffs p ��U  0��U  pjustforfun_justforfun_ ��U  0��U  ���U  p��U  0��U  ���i�  9! /       Meeting                        This_stuffs_This_stuffs_                                     D<�j�  (D /       Workout ffs ����U  P���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  K��j�  }D /       Workout ffs ���U  ����U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ڥ�j�  �G /       Birthday U  @_��U  P���U  �`Some_stuffs_Some_stuffs_ �U  �b��U  @c��U  �c��U  �d��U  �؏j�  �G /       Some_stuffs 0���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  ŉ�j�  �I /      Workout     ���U  ����U  P�Some_stuffs_Some_stuffs_ �U  @���U  ���U  ���U  ����U  ��,k�  �o /      Meeting     ���U  ж��U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��2k�  Pq /       Some_stuffs �<��U  �=��U   >Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �A��U  X��k�  � /       Birthday    ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  Bz�k�  � /       Appointment ����U  @���U  ��Some_stuffs_Some_stuffs_ �U  ����U  ����U  @���U  ����U  ���k�  �� /      Appointment 0E��U  �E��U  pFSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �J��U  ��@l�  �� /       Birthday    `���U  ����U  `�justforfun_justforfun_ ��U   ���U  ����U  `���U  ����U  t�Hl�  �� /      Some_stuffs p��U  0��U  0Some_stuffs_Some_stuffs_ �U   +��U  �+��U  �/��U  p0��U  �M�l�  t� /      Some_stuffs ����U  0���U  P
Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  X�l�  �� /       Workout     ���U  ���U  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ��l�  ,� /       Some_stuffs ���U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  1 �m�  � /       Workout     `k��U   l��U  �lThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �q��U  r	�m�  F /       Appointment ���U  Ѓ��U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  Ј��U  �Ԏm�  � /      Meeting     �r��U  �s��U  @tThis_stuffs_This_stuffs_ �U  �v��U  �w��U  x��U  �x��U   i
n�  �+ /       Meeting     ����U  P���U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  E�n�  l, /      Workout �U  0���U  ����U  �justforfun_justforfun_ ��U  p���U  ����U  p���U  0���U  �~#n�  2 /       Birthday    P���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �3)n�  �3 /       Birthday    ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  ����U  ����U  ����U  x#�n�  [X /       Some_stuffs �K��U  0L��U  �Ljustforfun_justforfun_ ��U  �O��U  pP��U  �P��U  �Q��U  �Go�  �| /       Workout     p��U  0��U  0This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p0��U  �&Vo�  �� /       Meeting     �O��U  pP��U  �PSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �U��U  ��]o�  r� /      Birthday    ���U  0 ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �3��U  K_�o�  ݠ /       Some_stuffs  ��U  ���U   justforfun_justforfun_ ��U   ��U  ���U   ��U  ���U  ���o�  k� /       Appointment ����U  ����U   �Some_stuffs_Some_stuffs_ �U  ����U   ���U  ����U  `���U  x��o�  �� /       Workout ent P���U  ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  ��o�  �� /      Appointment p��U  0��U  0This_stuffs_This_stuffs_ �U   +��U  �+��U  �/��U  p0��U  :op�  s� /       Some_stuffs ���U  p��U  0Some_stuffs_Some_stuffs_ �U  ���U  0 ��U  � ��U  p!��U  YH�p�  '� /       Workout      ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  p���U  ���U  ж��U  ��p�  '� /      Meeting �U  p��U  0��U  �This_stuffs_This_stuffs_ �U  ���U  ���U  p��U  ���U  �'�p�  +� /       Some_stuffs 0���U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �cq�  �� /       Meeting     л��U  ����U  ��This_stuffs_This_stuffs_ �U  0���U  ���U  ����U  p���U  |$q�  �� /       Birthday nt @��U  ���U  @This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ��U  �Zq�  � /       Workout �U  p���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  �}q�  �� /      Workout     ����U  ����U   �This_stuffs_This_stuffs_ �U  Ћ��U  ����U   ���U  ����U  A�#q�  �� /       Some_stuffs ��U  ���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0��U  7E�q�  " /      Meeting     @ ��U  � ��U  @!Some_stuffs_Some_stuffs_ �U  �#��U  �$��U   %��U  �%��U  +�q�  � /       Meeting     P��U  ���U  PSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p#��U  �q�  _ /       Meeting �U  �s��U   t��U  �tSome_stuffs_Some_stuffs_ �U  w��U  �w��U  x��U  �x��U  �u�q�  A /       Appointment ����U  @���U  �justforfun_justforfun_ ��U  P���U  ���U   ���U  ����U  ���q�   /       Some_stuffs ��	��U  `�	��U  ��	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   �	��U  ��>r�  (? /      Some_stuffs ���U  @	��U  �	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  )�Jr�  IB /       Meeting �U  ���U  ����U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ���r�  Qe /      Some_stuffs @���U   ���U  ��Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  A�hs�  h� /       Workout �U  E��U  �E��U  PFSome_stuffs_Some_stuffs_ �U  PH��U  I��U  �I��U  �J��U  *�is�  �� /       Workout �U  ����U  P���U  �justforfun_justforfun_ ��U  ����U  `���U  Э��U  P���U  {Iks�  � /       Meeting     p���U  0���U  ��Some_stuffs_Some_stuffs_ �U  ���U  ����U  ���U  ����U  $�os�  8� /      Meeting     p ��U  0��U  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0��U  �t�  #� /      Workout     0���U  ����U  ��justforfun_justforfun_ _ �U  0���U  ����U  p���U  ����U  Iћ��  �( /       Meeting     ����U  p���U  0�justforfun_justforfun_ ��U  ����U  0���U  ���U  ����U  �����  Z�( /      Meeting �U  ����U  0���U  ��This_stuffs_This_stuffs_ �U  ����U  p���U  0���U  ����U  �ݤ��  n�( /       Birthday    ���U  Ћ��U  ��This_stuffs_This_stuffs_ �U  Э��U  P���U   ���U  ����U  e����  @%) /      Workout     `��U   ��U  �Some_stuffs_Some_stuffs_ �U  0��U  ���U  p��U  ���U  x�Ƞ�  )) /       Appointment  ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  %[��  �N) /      Workout     ���U   ��U  �Some_stuffs_Some_stuffs_ �U   ��U  ���U   ��U  ���U  rp��  T) /       Birthday U  `���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  T��  �r) /      Meeting     ����U  `���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ����  �t) /       Workout �U   ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  Н��U  ����U  ����U  p���U  �#���  ,�) /       Workout     ���U  ����U  P�Some_stuffs_Some_stuffs_ �U  ���U  Ш��U  ����U  P���U  T	���  ��) /      Birthday U  0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  ���  ��) /       Some_stuffs 0f��U  �g��U  �ijustforfun_justforfun_ _ his_stuffs_This_stuffs_ �U  �t��U  ���  ��) /       Workout     ���U  о��U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  
�,��  ��) /       Some_stuffs p���U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  |B4��  ��) /      Birthday    �?��U  P@��U  ASome_stuffs_Some_stuffs_ �U  �C��U  �D��U  E��U  �E��U  C�6��  h�) /       Birthday    ����U  P���U  ��This_stuffs_This_stuffs_ �U  ���U  ����U  P���U  ����U  h����  �) /       Appointment ����U  P���U  �justforfun_justforfun_ ��U  P���U  ����U  ����U  P���U  1�H��  ~* /       Appointment @S��U  �S��U  @TThis_stuffs_This_stuffs_ �U  @V��U   W��U  �W��U  @X��U  *d��  �* /       Meeting     ����U  @���U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  se��  �* /       Workout     @���U   ���U  ��justforfun_justforfun_ ��U  ����U  @���U   ���U  ����U    k��  T* /       Birthday fs �}��U  `~��U   justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  `���U  �d��  �6* /       Meeting                        Some_stuffs_Some_stuffs_                                     ���  �6* /       Workout     @ ��U  � ��U  @!This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �%��U  `���  �6* /       Some_stuffs ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  @���U  0���U   ���U  �b��  e7* /       Birthday    p ��U  0��U  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0��U  ����  `;* /       Meeting     P��U  ��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0��U  �����  �;* /       Meeting     p���U  ����U  p�justforfun_justforfun_ ��U  ����U  0���U  ����U  ����U  !T���  =* /      Appointment ���U   ��U  �justforfun_justforfun_ ��U  �	��U  �
��U   ��U  ���U  9ꖥ�  d* /       Some_stuffs p���U  ����U  p�justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ����U  �x���  yd* /       Appointment  ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  Н��U  ����U  ����U  p���U  ����  ��* /       Workout     ���U  ����U  0�Some_stuffs_Some_stuffs_ �U   ���U  ����U  ����U  @���U  �U��  p�* /       Appointment �)��U  0*��U  �*Some_stuffs_Some_stuffs_ �U  p-��U  0.��U  �.��U  p/��U  h�(��  q�* /       Meeting �U   ���U  ����U  ��justforfun_justforfun_ ��U  Н��U  ����U  ����U  p���U  a����  ��* /       Some_stuffs E��U  �E��U  PFSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �J��U  N����  ��* /      Workout     0u��U  �u��U  pvThis_stuffs_This_stuffs_ �U  0y��U  �y��U  pz��U  0{��U  �C���  ��* /       Meeting �U  ���U  p��U  0This_stuffs_This_stuffs_ �U  0��U  ���U  0��U  ���U  a�P��  <�* /       Meeting     ���U  0��U  �This_stuffs_This_stuffs_ �U  ���U  ���U  p��U  0��U  �WU��  \�* /      Birthday    @���U  ����U  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  a����  ��* /       Workout     ����U  `���U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `���U  � ���  �+ /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �&w��  � + /       Some_stuffs `?��U   @��U  �Njustforfun_justforfun_ ��U  �B��U  pC��U  0D��U  �D��U  �ބ��  $+ /      Workout      ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ����  $+ /       Workout     P[��U  \��U  �`This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �h��U  ���  �J+ /      Appointment ����U  p���U  0�Some_stuffs_Some_stuffs_ �U  ���U  ����U  ����U  @���U  d����   n+ /      Meeting     0���U  ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  qs���  �q+ /       Appointment PH��U  I��U  �ISome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  �N��U  �@��  ��+ /       Meeting  fs е��U  ����U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  B�H��  ȗ+ /       Some_stuffs ����U  0���U  P
justforfun_justforfun_ ��U  ����U   ���U  ����U  @���U  ��P��  ڙ+ /       Some_stuffs 0���U   ���U  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  �xS��  }�+ /      Birthday                       justforfun_justforfun_                                       5pU��  ��+ /       Appointment �
��U  ���U  pSome_stuffs_Some_stuffs_ �U  ���U  ���U  p��U  0��U  4:^��  >�+ /       Some_stuffs @"��U   #��U  �#Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �'��U  n�^��  Q�+ /       Some_stuffs ����U  `���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �۪�  0�+ /       Workout      o��U  �o��U  �pjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  �u��U  ����  E�+ /      Workout     ����U  `���U  ��Some_stuffs_Some_stuffs_ �U  ���U  `��U  ��U  ���U  ��|��  ��+ /      Birthday    0���U  ����U  p�This_stuffs_This_stuffs_ �U  ����U  ����U  p���U  ����U  �ď��  v�+ /       Workout �U  ����U  @���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �_��  V
, /       Meeting     �Z��U  �[��U  @\This_stuffs_This_stuffs_ �U  `_��U   `��U  �`��U  `a��U  �u	��  �
, /      Workout ffs  ���U  ����U  ��Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  ж��U  �)��  �, /       Workout     �Z��U  �[��U  @\This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  �`��U  �栬�  b1, /       Appointment '	��U  �'	��U  (	Some_stuffs_Some_stuffs_ �U  �*	��U   +	��U  �+	��U   ,	��U  1ѡ��  �1, /       Meeting     ���U  p���U  0�This_stuffs_This_stuffs_ �U  ����U  p���U  ����U  p���U  ���  7, /      Some_stuffs ���U  0��U  �justforfun_justforfun_ _ �U  p��U  0��U  ���U  0��U   :��  �X, /       Some_stuffs `o��U   p��U  �pjustforfun_justforfun_ ��U  �s��U  pt��U  0u��U  �u��U  ��B��  �Z, /      Meeting ent ���U  ж��U  ��justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  ����U  CD��  ([, /       Some_stuffs ���U  0��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0��U  2iY��  �`, /       Appointment ���U  p��U  0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �!��U  ���  )�, /      Birthday    @���U  ����U  @�This_stuffs_This_stuffs_ �U  ����U   ���U  ����U  ����U  �o��  ��, /       Birthday    0���U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U   .s��  ��, /       Meeting     �
��U  ���U  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0��U  �i��  ��, /       Some_stuffs ����U  ���U  ��This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  @���U  �
��  ��, /      Some_stuffs �l��U  `m��U   justforfun_justforfun_ ��U  �p��U  �q��U  0r��U  �r��U  ��G��  � - /      Meeting     0���U  ����U  p�Some_stuffs_Some_stuffs_ �U  P
��U  �
��U  @���U  ����U  P4H��  � - /       Birthday    �/��U  p0��U  �4This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �F��U  �}L��  �!- /       Workout     p���U  ����U  ��This_stuffs_This_stuffs_ �U  0���U  ����U  ����U  0���U  �̰�  �B- /       Some_stuffs е��U  ����U  �Some_stuffs_Some_stuffs_ �U  ����U  ����U  ���U  ����U  ��հ�  E- /      Appointment @p��U   q��U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  v��U  ��w��  }n- /      Birthday    �G��U  0H��U  �Hjustforfun_justforfun_ ��U  �K��U  0L��U  �L��U  �M��U  z�!��  �8 /       Birthday fs ����U  ���U  ��justforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U  0���U  ;z5��  8 /       Birthday    @[��U  �[��U  `\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p`��U  �18��  �8 /       Workout     @���U  ����U  @�This_stuffs_This_stuffs_ �U  ����U  P���U  д��U  P���U  ��9��  :8 /      Workout     `���U   ���U  ��This_stuffs_This_stuffs_ �U  `���U   ���U  ����U   ���U  �Z���  �?8 /      Meeting     ����U  P���U  мThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  )#���  	@8 /       Some_stuffs ���U  `��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �#��U  a�_��  |j8 /       Birthday U  P�	��U  ��	��U  P�	This_stuffs_This_stuffs_ �U  ��	��U   �	��U  ��	��U   �	��U  P>b��  k8 /       Meeting     �z��U  `{��U   |This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  Z<���  ��8 /       Workout     p���U  0���U  �justforfun_justforfun_ ��U  P���U  ���U  Р��U  ����U  p����  ��8 /       Appointment ���U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  n���  C�8 /      Some_stuffs p��U  0��U  �Some_stuffs_Some_stuffs_ �U  0��U  ���U  ���U  p��U  ���  ��8 /       Some_stuffs p��U  0��U  �justforfun_justforfun_ ��U  ���U  0��U  ���U  p��U  5���  ¶8 /      Workout �U  @f��U  �f��U  @gjustforfun_justforfun_ ��U  �i��U  @j��U   k��U  �k��U  �I���  k�8 /       Birthday    P[��U  \��U  �`justforfun_justforfun_ ��U   l��U  �l��U  �g��U  �h��U  �)���  o�8 /       Meeting      ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  [���  '�8 /       Workout     �1��U   2��U  �2This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P7��U  ]a"��  ��8 /      Birthday U  PO��U  �O��U  �PSome_stuffs_Some_stuffs_ �U  �R��U  PS��U  T��U  �T��U  b9��  ��8 /       Meeting ffs  ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  X�9��  ��8 /       Appointment �L��U  �M��U  @^justforfun_justforfun_ ��U  �P��U  �Q��U  pR��U  �R��U  ܺV��  �,9 /      Some_stuffs ����U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��k��  #29 /       Some_stuffs �t��U  �u��U  vjustforfun_justforfun_ ��U  `y��U   z��U  �z��U  `{��U  ����  /R9 /       Appointment �z��U  `{��U   |Some_stuffs_Some_stuffs_ �U  p��U  0���U  ����U  ����U  �����  �W9 /      Meeting �U  p���U  0���U  ��This_stuffs_This_stuffs_ �U  P���U  ���U  ����U  P���U  z����  �W9 /       Birthday    `���U  ���U  ��This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ���U  Ǆ��  z9 /      Birthday    00��U  �0��U  p1Some_stuffs_Some_stuffs_ �U  04��U  �4��U  05��U  �5��U  P����  �}9 /       Birthday    P-��U  �-��U  �.This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �2��U  T� ��  ��9 /      Some_stuffs  E��U  �F��U  0KThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  \��U  �y"��  m�9 /       Birthday    pB��U  �B��U  �CThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �G��U  `���  �9 /       Meeting      2��U  �2��U   3Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   7��U  �JV��  :�9 /       Workout     ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  �sb��  W�9 /       Workout     0y��U  �y��U  pzSome_stuffs_Some_stuffs_ �U  �|��U  �}��U  0~��U  ����U  4����  �: /      Birthday                       justforfun_justforfun_                                       �[���  �: /       Meeting     �g��U  �h��U  pjSome_stuffs_Some_stuffs_ �U  �m��U  @n��U   o��U  �o��U  4����  b?: /      Appointment ����U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �r���  eA: /       Birthday    �z��U  `{��U   |This_stuffs_This_stuffs_ �U  p��U  0���U  ����U  ����U  �w��  �c: /      Workout                        This_stuffs_This_stuffs_                                     ��$��  �g: /       Some_stuffs  ��U  ���U   justforfun_justforfun_ _ �U   ��U  ���U   ��U  ���U  �&��  �g: /       Workout     ����U  ����U   �Some_stuffs_Some_stuffs_ �U  Ћ��U  ����U   ���U  ����U  +�*��  )i: /       Workout     ����U  P���U  ��Some_stuffs_Some_stuffs_ �U  ���U  ����U  ���U  ����U  @����  h�: /       Workout     Ц��U  ����U  �Some_stuffs_Some_stuffs_ �U  Ъ��U  ����U  P���U  ���U  �����  ��: /      Meeting     �f	��U  `g	��U  �g	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �k	��U  fF��  ı: /      Birthday    �
��U  ���U  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0��U  P���  r�: /       Appointment `���U   ���U  ��Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   ���U  �kw��  ��: /      Workout     ����U  P���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  PȌ��  R; /       Workout �U  p���U  ���U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  
Q
��  u%; /       Workout     ���U  p��U  0This_stuffs_This_stuffs_ �U  ���U  p��U  0��U  ���U  �>��  �*; /       Birthday    ����U  `���U   �justforfun_justforfun_ ��U  `���U   ���U  ����U  ����U  55,��  ".; /      Workout     е��U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ���  �S; /      Meeting     �(��U  P)��U  �)This_stuffs_This_stuffs_ �U  �+��U  �,��U   -��U  �-��U  @����  hT; /       Workout     Н��U  ����U  ��This_stuffs_This_stuffs_ �U  p���U  0���U  ���U  ����U  D+C��  �u; /      Some_stuffs                    justforfun_justforfun_                                       acD��  �u; /       Workout     ���U  ����U  P�This_stuffs_This_stuffs_ �U  @���U  ���U  ���U  ����U  �I��  w; /       Workout     ����U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  p���U  0���U  ����U  �*R��  cy; /       Meeting ent p���U  0���U  ��justforfun_justforfun_ _ �U  p���U  ����U  ����U  0���U  �c���  ��; /       Birthday    ����U  @���U  ��This_stuffs_This_stuffs_ �U   ���U  ����U  @ ��U  � ��U  t���  Y�; /      Workout     @^��U  �^��U  �OThis_stuffs_This_stuffs_ �U  pR��U  �R��U  �S��U  pT��U  )j���  i�; /       Workout ffs ����U  p���U  �justforfun_justforfun_ _ �U  ���U  ����U  @���U  ����U  ��m��  �; /      Appointment P��U  ���U  PSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p#��U  �v��  �; /       Some_stuffs  ���U  ����U  @�justforfun_justforfun_ ��U  ����U   ���U  ����U  @���U  �|��  ��; /       Appointment �
��U  ���U  pThis_stuffs_This_stuffs_ �U  ���U  ���U  p��U  0��U  ����  k�; /       Workout     ���U  ����U  P�justforfun_justforfun_ ��U  ���U  ����U  ����U  P���U  �,��  ��; /       Birthday nt ��U  ���U  This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P��U  �"��  %�; /       Birthday U  ���U   ��U  �This_stuffs_This_stuffs_ �U   ��U  ���U  0��U  ���U  ��(��  ��; /       Meeting      &��U  �&��U  0justforfun_justforfun_ _ �U  0��U  ���U  p��U  ���U  lf���  �< /      Appointment p ��U  0��U  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0��U  ᧴��  �< /       Workout ffs `y��U   z��U  �zThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  0���U  �`x��  P�< /      Appointment е��U  ����U  �This_stuffs_This_stuffs_ �U  ����U  ����U  ���U  ����U  ���  �[G /       Some_stuffs K��U  �K��U  PLThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Q��U  ����  X^G /       Birthday    x��U  �x��U  �yjustforfun_justforfun_ ��U  |��U  �|��U  �}��U  ~��U  .���  �`G /      Meeting     P���U  ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  e�S�  ��G /       Meeting     �2��U   3��U   4This_stuffs_This_stuffs_ �U  `6��U   7��U  �7��U  `8��U  �T�  .�G /      Birthday    ����U  @���U   �This_stuffs_This_stuffs_ �U  @���U  ����U  @���U  ����U  4'Y�  ^�G /       Birthday fs 0��U  ���U  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �"��U  Y�\�  G�G /       Meeting     ����U  p���U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0��U  ;�g�  �G /       Birthday    ����U  `���U  ЭThis_stuffs_This_stuffs_ �U  `���U  ����U  `���U  ����U  �m�  ��G /       Birthday    p ��U  0��U  pjustforfun_justforfun_ ��U  0��U  ���U  p��U  0��U  0��  ~�G /       Birthday    ����U  P���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  pݢ�  ��G /       Birthday    ����U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  ���  ��G /      Appointment �Z��U  �[��U  @\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �`��U  y#�  ��G /       Workout      k��U  �k��U  �lSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   q��U  �:1�  8�G /       Meeting     �v��U  �w��U  xjustforfun_justforfun_ ��U  �z��U  P{��U  |��U  �|��U  L���  �H /      Appointment 0���U   ���U  @�This_stuffs_This_stuffs_ �U  p���U  0���U  ����U  `���U  �=��  �!H /       Meeting     @���U   ���U  ��Some_stuffs_Some_stuffs_ �U  0���U  ����U  P���U  ���U  �V]�  IH /       Some_stuffs 0��U  ���U  �justforfun_justforfun_ ��U  ���U  p��U  0��U  ���U  �ic�  �JH /      Some_stuffs @\��U   ]��U  �]This_stuffs_This_stuffs_ �U  �`��U  `a��U   b��U  �b��U  pg��  rH /       Appointment ����U  ����U   �This_stuffs_This_stuffs_ �U  @���U  ����U  ����U   ���U  �҈�  ��H /       Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             Ka��  �H /       Appointment �L��U  �M��U  @NSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   R��U  ]���  K�H /      Meeting      ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ж��U  ���  O�H /       Workout     ���U  @���U  �Some_stuffs_Some_stuffs_ �U  @���U  ���U  p���U  ���U  ��"�  #�H /       Some_stuffs P���U  ����U  ��This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  P���U  �\'�  M�H /       Some_stuffs �N��U  PO��U  0ASome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �E��U  ݁*�  �H /      Some_stuffs ����U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  ,p6�  )�H /       Workout     ����U  `���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ;9�  ��H /       Meeting     ���U  p���U  0�Some_stuffs_Some_stuffs_ �U  p���U  ���U  ����U  p���U  +��  ��H /      Birthday    @\��U   ]��U  �]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �b��U  A���  h�H /       Appointment ���U  ����U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  �1��  D�H /       Birthday    E��U  �E��U  PFThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �J��U  "�J�  �I /       Birthday    �	��U  0
��U  �
justforfun_justforfun_ ��U  ���U  0��U  ���U  ���U  lP�  Y
I /      Birthday                       Some_stuffs_Some_stuffs_                                     �0R�  �
I /       Meeting     @���U  ����U  @�Some_stuffs_Some_stuffs_ �U  ����U  P���U  д��U  P���U  �i^�  �I /       Meeting     `V��U   W��U  �WSome_stuffs_Some_stuffs_ �U  �Z��U  �[��U  @\��U   ]��U  �^��  �4I /      Workout     pF��U  0G��U  �GThis_stuffs_This_stuffs_ �U  0J��U  �J��U  �K��U  0L��U  (r}�  iWI /       Meeting      1��U  �1��U  �2This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   7��U  uj�  �WI /      Meeting     ���U  й��U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  l��  1~I /       Appointment 0���U  ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  b�#�  ��I /       Appointment 0���U  ����U  p�Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   ���U  �<*�  ��I /       Birthday U  @���U   ���U  ��This_stuffs_This_stuffs_ �U  ����U  @���U   ���U  ����U  �+�  ڃI /       Meeting �U  ����U  0���U  ��justforfun_justforfun_ ��U  ����U  ����U  ���U  ����U  -&3�  �I /      Some_stuffs  E��U  �F��U  0Kjustforfun_justforfun_ ��U  �U��U  �V��U  P[��U  \��U  ~��  ?�I /       Appointment ����U  P���U  �justforfun_justforfun_ ��U  P���U  ����U  ����U  P���U  �o��  שI /       Appointment p ��U  0��U  pjustforfun_justforfun_ ��U  0��U  ���U  p��U  0��U  N���  A�I /      Workout     @���U  ����U  ��Some_stuffs_Some_stuffs_ �U   ���U  ����U  @ ��U   ��U  ��K �  ��I /       Some_stuffs @���U  ����U  ��Some_stuffs_Some_stuffs_ �U   ���U  ����U  @ ��U   ��U  �zQ �  :�I /      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��Y �  Y�I /       Some_stuffs p ��U  0��U  pThis_stuffs_This_stuffs_ �U  0��U  ���U  p��U  0��U  ��� �  =�I /      Birthday    0���U   ���U  @�justforfun_justforfun_ ��U  p���U  0���U  ����U  `���U  I�w!�  �J /       Workout     p���U  0���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  h݈!�  �J /       Appointment  ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  `���U   ���U  ����U  �k�!�  �J /      Appointment 0���U  ����U  p�Some_stuffs_Some_stuffs_ �U  ���U  ����U  0���U  ����U  ��"�  �@J /       Appointment ���U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �!"�  $FJ /      Some_stuffs ��U  ���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0��U  �""�  -FJ /       Workout     p��U  0��U  0This_stuffs_This_stuffs_ �U   +��U  �+��U  �/��U  p0��U  �"�  �gJ /       Meeting ent ����U  `���U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `���U  j��"�  �oJ /       Workout     ����U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  9;�"�  �pJ /       Birthday    0���U  ����U  ��This_stuffs_This_stuffs_ �U  p���U  0���U  ����U  p���U  ��A#�  ׏J /       Some_stuffs ���U  p���U  �justforfun_justforfun_ ��U  p���U  ���U  p���U   ���U  J>K#�  =�J /       Meeting     ����U  @���U   �Some_stuffs_Some_stuffs_ �U   ���U  p���U  ����U  `���U  Xd`#�  ��J /       Meeting     0���U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �b�#�  <�J /      Appointment  ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  �$�  �J /      Appointment ����U  @���U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  �%�  $K /       Some_stuffs �,��U  �-��U  @.Some_stuffs_Some_stuffs_ �U   1��U  �1��U  �2��U   3��U  �P�%�  �-K /      Appointment �z��U  P{��U  |This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  �c�%�  �-K /       Appointment 0f��U  �g��U  �iSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  �t��U  ��%�  �1K /       Appointment ����U  ����U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  +O>&�  �SK /       Appointment Н��U  p���U  0�Some_stuffs_Some_stuffs_ �U  ����U  p���U  0���U  ���U  H�>&�  �SK /       Workout �U   ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  p���U  ���U  ж��U  ��H&�  CVK /       Appointment ����U  `���U  @�Some_stuffs_Some_stuffs_ �U  ����U  ����U  ����U  `���U  e�R&�  �XK /      Meeting      o��U  �o��U  �pjustforfun_justforfun_ ��U  Ps��U  t��U  �t��U  �u��U  ҅�&�  �zK /       Workout ent �(��U  �)��U  @*Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �.��U  y��&�  ~K /       Some_stuffs ����U  ����U  0�Some_stuffs_Some_stuffs_ �U  `���U  �.	��U  `���U  ���U  ��&�  C�K /       Workout     �N��U  PO��U  0ASome_stuffs_Some_stuffs_ �U  0D��U  �D��U  0E��U  �E��U  0�o'�  ��K /       Some_stuffs  ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  p���U  ���U  ж��U  ��s'�  ͢K /       Birthday     ���U  ����U  `�Some_stuffs_Some_stuffs_ �U  `���U   ���U  ����U   ���U  �}'�  N�K /      Meeting     ���U  й��U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  cf'�  ��K /       Meeting ent �	��U  �
��U   Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  N(�  ?�K /       Appointment P[��U  \��U  �`Some_stuffs_Some_stuffs_ �U   l��U  �l��U  �g��U  �h��U  �h(�  ��K /      Meeting     ���U  ����U  0�Some_stuffs_Some_stuffs_ �U   ���U  ����U  ����U  @���U  (�  x�K /       Workout     ����U  0���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  |ۦ(�  _�K /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �*TR�  ��V /       Workout     ���U  о��U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ЛrR�  ��V /       Some_stuffs p���U  0���U  ��This_stuffs_This_stuffs_ �U  0���U  ���U  ����U  p���U   ��R�  ��V /       Workout     0���U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  ��R�  /�V /       Some_stuffs PG��U  �G��U  PHSome_stuffs_Some_stuffs_ �U  K��U  �K��U  PL��U  M��U  �ˑS�  �V /      Birthday     +��U  �+��U  �/Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �?��U  9�S�  ��V /       Birthday nt  >��U  �>��U  `?Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  pC��U   g�T�  �9W /       Some_stuffs ����U  P���U  ��Some_stuffs_Some_stuffs_ �U  P���U  ����U  P���U  ����U  i�T�  J=W /       Appointment е��U  ����U  �This_stuffs_This_stuffs_ �U  ����U  ����U  ���U  ����U  �pU�  xhW /       Workout     ����U  p���U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  ��U�  όW /       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �V�  ^�W /      Workout     @X��U  �X��U  �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ^��U  (��V�  ɯW /       Workout �U  0f��U  �g��U  �iSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �t��U  :��V�  S�W /       Appointment �;��U  `<��U  �<justforfun_justforfun_ ��U  `?��U   @��U  �N��U  PO��U  �ʐV�  a�W /       Meeting     ����U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  @���U   ���U  ����U  cE W�  �W /       Workout     0p��U  �p��U  pqThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Pu��U  �b,W�  6�W /       Meeting     ����U  `���U  ЭSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��,W�  Z�W /      Birthday     ���U  ����U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  ��2W�  ��W /       Some_stuffs `V��U   W��U  �WThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ]��U  Y�2W�  ��W /       Appointment �%��U  0&��U  �&Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p+��U  �=<W�  E�W /       Some_stuffs �i��U  @j��U   kSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �o��U  ��W�  �W /       Birthday     ���U  ����U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  м��U  `[�W�  � X /       Appointment 0f��U  �g��U  �ijustforfun_justforfun_ ��U  �p��U  �q��U  �s��U  �t��U  R��X�  rJX /       Some_stuffs ����U   ���U  ��justforfun_justforfun_ _ his_stuffs_This_stuffs_ �U  @��U  ���X�  �LX /       Workout     ����U  `���U   �justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ����U   ?�X�  `MX /       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             յ�X�  �NX /      Workout ent ����U  @���U  �justforfun_justforfun_ ��U  P���U  ���U   ���U  ����U  Ln�X�  =PX /       Some_stuffs @'��U  �'��U  @(Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �,��U  ��Y�  5vX /       Workout     `:��U   ;��U  �;This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   @��U  ��Z�  �X /       Some_stuffs                    Some_stuffs_Some_stuffs_                                     �Z�  Y�X /      Appointment p��U  0��U   &This_stuffs_This_stuffs_ �U  ���U  p��U  0��U  ���U  C˻Z�  ��X /       Some_stuffs �+��U   ,��U  �,This_stuffs_This_stuffs_ �U  �/��U  @0��U   1��U  �1��U  �.�Z�  ��X /       Meeting �U   ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  `���U   ���U  ����U  9[�Z�  ��X /       Birthday    p���U  ����U  ��Some_stuffs_Some_stuffs_ �U  p���U  ����U  p���U  ����U  v�Z�  ��X /      Workout     0"��U  �<��U  0$This_stuffs_This_stuffs_ �U  �&��U  �'��U  0(��U  �(��U  (N[�   �X /       Workout     �W��U  �X��U  @YThis_stuffs_This_stuffs_ �U  @\��U   ]��U  �]��U  �n��U  ��X[�  ��X /       Meeting      ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  `���U  ����U  `���U  �X`[�  ��X /      Workout     ����U   ���U  ��This_stuffs_This_stuffs_ �U  ����U  p���U  0���U  ���U  ��[�  LY /       Workout     �6��U   7��U  �7justforfun_justforfun_ ��U  P9��U  �9��U  p:��U  0;��U  t��[�  �Y /      Birthday U  ����U  ����U  ��justforfun_justforfun_ ��U  ����U  p���U  0���U  ����U  �!�\�  �7Y /       Appointment ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  ܷ�\�  �<Y /      Appointment ��U  ���U  �Some_stuffs_Some_stuffs_ �U  ���U  ���U  p��U  0��U  �Z(]�  ebY /      Meeting �U  �B��U  pC��U  0DSome_stuffs_Some_stuffs_ �U  pF��U  0G��U  �G��U  0H��U  �,�]�  $�Y /       Workout     ����U  P���U  ��Some_stuffs_Some_stuffs_ �U  P���U  ����U  P���U  ����U  �Ʊ]�  ��Y /      Birthday    `y��U   z��U  �zSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  0���U  @��]�  (�Y /       Birthday    �z��U  `{��U   |This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �,�]�  x�Y /       Workout     0���U  ���U  ��justforfun_justforfun_ ��U  ���U  p���U  0���U  ����U  ���]�  %�Y /       Birthday    �(��U  P)��U  �)Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �-��U  ��?^�  ��Y /       Appointment ����U  @���U  P�Some_stuffs_Some_stuffs_ �U  P���U  Т��U  ����U  P���U  ��@^�  ;�Y /      Some_stuffs ����U  p���U  0�justforfun_justforfun_ ��U  0���U  ����U  p���U  0���U  j
L^�  �Y /       Appointment 0��U  ���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0 ��U  ��^�  2�Y /      Appointment �t��U  �u��U  vThis_stuffs_This_stuffs_ �U  `y��U   z��U  �z��U  `{��U  �xx_�  ��Y /       Birthday    @���U  ����U  @�This_stuffs_This_stuffs_ �U  ����U  P���U  д��U  P���U  ��~_�  ��Y /       Workout     ����U  0���U  ��Some_stuffs_Some_stuffs_ �U  ����U  0���U  ����U  ����U  N�_�  ��Y /       Some_stuffs ���U  ���U   This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ��U  �m�_�  ��Y /      Meeting      ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  Į`�  �"Z /      Birthday     ���U  ����U  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  �ڦ`�  cGZ /       Appointment �p��U   q��U  �wThis_stuffs_This_stuffs_ �U  �t��U  �u��U  v��U  �v��U  ���`�  %KZ /      Birthday fs 0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  2ظ`�  �KZ /       Workout     ����U  @���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  a5�`�  MZ /       Workout     ����U  p���U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �v�`�  �NZ /       Appointment ����U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  ��:a�  LmZ /       Birthday     ���U  ����U   �Some_stuffs_Some_stuffs_ �U  ����U  p���U  Љ��U  ����U  �!Xa�  �tZ /       Appointment ����U  p���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  �]a�  .vZ /      Birthday    ���U  ����U  `�justforfun_justforfun_ ��U  ����U  @���U   ���U  ����U  ���a�  ��Z /      Workout     @��U  ���U  @Some_stuffs_Some_stuffs_ �U   ��U  ���U   	��U  �	��U  H��a�  ��Z /       Birthday U  P[��U  \��U  �`This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �h��U  ��zb�  /�Z /       Workout     @���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  ���b�  E�Z /      Birthday    ���U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  �A�b�  k�Z /       Meeting      ��U  ���U   This_stuffs_This_stuffs_ �U  @��U  ���U  @��U  ���U  �_c�  ��Z /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             1&c�  ��Z /       Workout     ����U  @���U  �Some_stuffs_Some_stuffs_ �U  P���U  ���U   ���U  ����U  
J�c�  [ /       Some_stuffs 0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  ֧c�  ?[ /       Workout     p"��U  �"��U  �#This_stuffs_This_stuffs_ �U  @'��U   (��U  �(��U  �)��U  `òc�  [ /      Birthday U  0��U  ���U  �This_stuffs_This_stuffs_ �U  0"��U  �<��U  0$��U  �$��U  8еc�  �[ /       Some_stuffs p���U  0���U  ��justforfun_justforfun_ ��U  ����U  ����U   ���U  ����U  Ҷc�  [ /       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �V�c�  7[ /       Appointment  o��U  �o��U  �pSome_stuffs_Some_stuffs_ �U  Ps��U  t��U  �t��U  �u��U  Đ��  ��e /      Appointment 0���U  ���U  ��justforfun_justforfun_ ��U  ����U  0���U  ���U  p���U  �����  �f /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ٶ���  7f /       Birthday    ���U  ����U  ��justforfun_justforfun_ ��U  0���U  ����U  ����U  p���U  ��!��  �-f /      Birthday fs ���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  (A��  �5f /       Some_stuffs @p��U   q��U   �justforfun_justforfun_ ��U  @t��U  �t��U  �u��U  v��U  ��B��  �5f /       Some_stuffs  9��U  �9��U  `:This_stuffs_This_stuffs_ �U  �<��U  �=��U   >��U  �>��U  �ݹ��  rTf /      Some_stuffs  ���U  ����U  ��This_stuffs_This_stuffs_ �U  0���U  ����U  ����U  p���U  i[Ώ�  �Yf /       Workout     ����U  ����U  P�Some_stuffs_Some_stuffs_ �U  ���U  ����U  ����U  P���U  �R��  �{f /       Appointment ����U  p���U  0�Some_stuffs_Some_stuffs_ �U  ����U  0���U  ����U  ����U  �Y��  3}f /      Meeting ffs ����U  ����U  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  ����  ȣf /      Appointment p��U  0��U  0justforfun_justforfun_ ��U   +��U  �+��U  �/��U  p0��U  0n���  ��f /       Appointment                    Some_stuffs_Some_stuffs_                                     ᵆ��  l�f /       Appointment 04��U  �4��U  05justforfun_justforfun_ ��U  p7��U  08��U  �8��U  p9��U  `G���  \�f /       Workout �U  p ��U  0��U  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0��U  �i+��  ��f /       Birthday nt ����U  P���U  дSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  p�2��  ��f /       Workout     �h��U   i��U  �iSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @n��U  =y���  wg /      Appointment P���U  ���U  p�Some_stuffs_Some_stuffs_ �U  ����U  ����U  @���U    ��U  hɒ�  �g /       Birthday nt pF��U  0G��U  �GThis_stuffs_This_stuffs_ �U  0J��U  �J��U  �K��U  0L��U  �>Ӓ�  �g /       Some_stuffs @��U   ��U  �justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ���U  ,�P��  �?g /      Meeting �U  @S��U  �S��U  @TThis_stuffs_This_stuffs_ �U  @V��U   W��U  �W��U  @X��U  QFR��  @g /       Some_stuffs 0��U  ���U  pjustforfun_justforfun_ ��U  ���U  ���U  0��U  ���U  ;]��  �Bg /       Appointment ����U  ����U  �justforfun_justforfun_ ��U  ����U  ����U  @���U  ����U  ���  0gg /       Meeting     �J��U  pK��U  �KThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �O��U  @Y��  Hhg /       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ]���  �kg /      Workout     `?��U   @��U  �NSome_stuffs_Some_stuffs_ �U  �B��U  pC��U  0D��U  �D��U  �q���  D�g /       Meeting �U  �}��U  `~��U   This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  �$���  x�g /       Workout �U  �)��U  0*��U  �*Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p/��U  n����  Ւg /      Appointment ���U  ����U  �This_stuffs_This_stuffs_ �U  P���U  ����U  P���U  ����U  �ѕ�  ��g /      Appointment P[��U  \��U  �`This_stuffs_This_stuffs_ �U   l��U  �l��U  �g��U  �h��U  ��\��  Xh /       Some_stuffs ����U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  @���U   ���U  ����U  ��e��  �	h /      Meeting �U  0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  Q���  �)h /       Some_stuffs ����U  p���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  ����  D-h /       Appointment 0���U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �~���  ;/h /      Meeting     pF��U  0G��U  �GSome_stuffs_Some_stuffs_ �U  0J��U  �J��U  �K��U  0L��U  �!z��  kPh /       Workout                        justforfun_justforfun_                                       >����  7Th /      Workout ent  ���U  ����U   �This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  ٴ���  �Vh /       Workout     ����U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ���  Mwh /       Meeting                        Some_stuffs_Some_stuffs_                                     ���  Zyh /       Appointment P���U  ���U  ��Some_stuffs_Some_stuffs_ �U  ���U  о��U  ����U  P���U  ����  �zh /      Birthday    �/��U  p0��U  �4Some_stuffs_Some_stuffs_ �U  �>��U  �?��U   E��U  �F��U  ?Ѳ��  w�h /      Some_stuffs �z��U  �{��U   |justforfun_justforfun_ ��U   ��U  ���U  `���U   ���U  Q����  ��h /       Birthday    ����U  `���U   �This_stuffs_This_stuffs_ �U  `���U   ���U  ����U  ����U  p
Ș�  �h /       Appointment ���U  p��U  0Some_stuffs_Some_stuffs_ �U  ���U  0 ��U  � ��U  �!��U  ro̘�  �h /       Meeting      ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  T�A��  �h /      Birthday    �)��U  0*��U  �*Some_stuffs_Some_stuffs_ �U  p-��U  0.��U  �.��U  p/��U  �ߙ�  v�h /       Birthday U   ���U  ����U  @ justforfun_justforfun_ ��U  ��U  ���U  ��U  ���U  :q��  s�h /       Birthday    @(��U  �(��U  p)This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �-��U  [6��  ��h /       Appointment ����U  ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  ��  `�h /       Birthday    p���U  ���U  ��This_stuffs_This_stuffs_ �U  0���U  ����U  ����U  0���U  �s��  ;i /      Workout     p���U  ����U  ��This_stuffs_This_stuffs_ �U  p���U  ����U  p���U  ����U  ��u��  �i /       Birthday    P[��U  \��U  �`Some_stuffs_Some_stuffs_ �U   l��U  �l��U  �g��U  �h��U  ����  yi /       Appointment ����U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ���  `?i /       Workout     ����U  `���U   �This_stuffs_This_stuffs_ �U  ����U  ����U   ���U  ����U  j�#��  q@i /       Meeting      >��U  �>��U  `?justforfun_justforfun_ ��U  0A��U  �A��U  �B��U  pC��U  ,*��  Bi /      Appointment p��U  0��U  �This_stuffs_This_stuffs_ �U  ���U  ���U  p��U  ���U  }r���  �ei /      Meeting     p��U  ���U  pThis_stuffs_This_stuffs_ �U  0��U  ���U  ���U  p��U  Hɺ��  gi /       Appointment ����U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  L���  �gi /       Workout     �Z��U  �[��U  @\This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  `a��U  ,�>��  �i /       Some_stuffs @t��U  �t��U  �uThis_stuffs_This_stuffs_ �U  x��U  �x��U  �y��U  Pz��U  )3C��  	�i /       Birthday nt  ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �W��  "�i /       Birthday nt ����U  @���U  ��justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ����U   �\��  ��i /       Meeting     �q��U  �r��U  �mjustforfun_justforfun_ ��U  �p��U   q��U  �w��U  �x��U  �7]��  ��i /      Appointment �f��U  �g��U  `hSome_stuffs_Some_stuffs_ �U  `k��U   l��U  �l��U  `m��U  ���  �i /       Birthday nt �K��U  pL��U   MSome_stuffs_Some_stuffs_ �U   O��U  �O��U   P��U  �P��U  t���  j�i /      Some_stuffs �,��U  �-��U  @.Some_stuffs_Some_stuffs_ �U   1��U  �1��U  �2��U   3��U  9ox��  3�i /       Appointment `���U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  �Q���  D�i /       Appointment `��U   ��U  �justforfun_justforfun_ ��U  0��U  ���U  p��U  ���U  ތ��  n�i /      Birthday    ���U  p��U  0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �!��U  M��  A�i /      Workout     pF��U  0G��U  �GSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0L��U   ���  tj /       Workout     �
��U  ���U  pThis_stuffs_This_stuffs_ �U  ���U  ���U  p��U  0��U  $i���  �$j /      Workout ffs ���U  ����U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �ݾ��  �,j /       Some_stuffs ���U  �	��U  �"Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  1�B��  ~Nj /       Birthday nt Н��U  ����U  ��This_stuffs_This_stuffs_ �U  p���U  0���U  ���U  ����U  �E��  EOj /      Appointment ���U  ����U  0�Some_stuffs_Some_stuffs_ �U   ���U  ����U  ����U  @���U  ����  �wj /       Some_stuffs 0���U  ����U  0�Some_stuffs_Some_stuffs_ �U  0���U  ����U  p���U  ����U  �.��  �yj /      Appointment ����U  `���U  ��Some_stuffs_Some_stuffs_ �U  ����U  `���U  е��U  ����U  �X���  �"u /      Birthday    p ��U  0��U  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0��U  /�#��  �Hu /      Some_stuffs ����U  ����U  ��This_stuffs_This_stuffs_ �U  ���U  ����U   ���U  ����U  _0��  �Ku /       Appointment ����U  0���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  :�4��  �Lu /       Appointment  R��U  �R��U  @SThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   W��U  Q�;��  �Nu /       Some_stuffs `���U   ���U  ��justforfun_justforfun_ ��U  `���U  ����U  `���U   ���U  �����  �ou /      Some_stuffs  ���U  ����U  �rjustforfun_justforfun_ ��U  �u��U  v��U  �v��U  �w��U  ҽ��  pu /       Meeting     �R��U  PS��U  TSome_stuffs_Some_stuffs_ �U  �q��U  `r��U   W��U  �W��U  1����  �tu /       Workout     ����U  @���U  ��Some_stuffs_Some_stuffs_ �U  ����U  @���U   ���U  ����U  ��Z��  O�u /      Meeting     `���U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  z#[��  [�u /       Some_stuffs �b��U  @c��U  �cjustforfun_justforfun_ ��U  �f��U  pg��U  0h��U  �h��U  9]a��  �u /       Workout      E��U  �F��U  0KThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  \��U  -3���  �u /      Some_stuffs �t��U  �u��U  vThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `{��U  (���  ��u /       Some_stuffs ����U  ����U  p�justforfun_justforfun_ ��U  ����U  @���U  ����U  ����U  �:���  :�u /      Birthday    p��U  0��U  �justforfun_justforfun_ ��U  ���U  ���U  p��U  ���U  ��"��  v /       Appointment 0���U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  H����  �5v /       Appointment е��U  ����U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  up���  �7v /      Appointment `5��U  �5��U  `6This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ;��U  B\���  (8v /       Workout     ���U  p��U  0Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  �!��U  e�U��  �[v /      Birthday U  �]��U  �n��U  `_Some_stuffs_Some_stuffs_ �U   b��U  �b��U   c��U  �c��U  h�c��  1_v /       Appointment ���U  ����U  `�Some_stuffs_Some_stuffs_ �U  ����U  @���U   ���U  ����U  D:���  �v /      Appointment 0r��U  �r��U  �sSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  px��U  tB���  �v /      Workout      ���U  ����U  `�Some_stuffs_Some_stuffs_ �U   ���U  ����U  `���U   ���U  �.2��  ��v /       Workout     ���U  @��U   Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  ����  1�v /      Some_stuffs �%��U  0&��U  �&This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p+��U  ��L��  �w /       Some_stuffs @\��U   ]��U  �]This_stuffs_This_stuffs_ �U  �`��U  `a��U   b��U  �b��U  pAN��  Fw /       Workout     0��U  ���U  pSome_stuffs_Some_stuffs_ �U  ���U  ���U  0��U  ���U  �E���  lDw /       Workout     �z��U  `{��U   |This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  g���  
Hw /       Meeting     p���U  ����U  ��This_stuffs_This_stuffs_ �U  p���U  ����U  p���U  ����U  D����  ,Kw /      Appointment ����U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �	���  �nw /      Some_stuffs                    justforfun_justforfun_                                       ��#��  x�w /       Workout     �R��U  PS��U  TSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �W��U  	(��  ��w /       Meeting     ����U  p���U  0�This_stuffs_This_stuffs_ �U  ����U  p���U  0���U  ����U  �c.��  0�w /      Appointment  ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  f���  C�w /      Birthday                       justforfun_justforfun_                                       Y���  '�w /       Birthday    @*��U   +��U  �+This_stuffs_This_stuffs_ �U  @.��U  �.��U  �/��U  @0��U  (pK��  )�w /       Meeting  nt p���U  ���U  p�Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  @���U  �����  0x /       Meeting     �{��U  0|��U  �|justforfun_justforfun_ _ his_stuffs_This_stuffs_ �U   ���U  �����  �x /       Appointment  l��U  �l��U  �gThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @n��U  ,�|��  M0x /      Workout �U  ����U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  ZG���  �3x /       Birthday    ����U  P���U  �justforfun_justforfun_ ��U  P���U  ����U  ����U  P���U  �2���  �5x /       Workout     �9��U  �:��U  p;Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P@��U  ؖ��   7x /       Appointment ���U  @��U  �Some_stuffs_Some_stuffs_ �U   ��U  ���U   ��U  ���U  �s)��  �\x /      Appointment @f��U  �f��U  @gjustforfun_justforfun_ _ �U  �i��U  @j��U   k��U  �k��U  X?1��  �^x /       Birthday                       This_stuffs_This_stuffs_                                     t{���  �|x /      Appointment ����U  @���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �����  �|x /       Meeting     P���U  ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  )���  ��x /       Some_stuffs ����U  P���U  ��justforfun_justforfun_ ��U  ���U  ����U  ���U  ����U  ��>��  ��x /       Workout     0���U   ���U  @�justforfun_justforfun_ ��U  p���U  0���U  ����U  `���U  �@��  
�x /       Birthday     P��U  �P��U   QSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �T��U  
�F��  ��x /       Some_stuffs 0���U  ����U  0�This_stuffs_This_stuffs_ �U  0���U  ����U  p���U  0���U  3�G��  ޥx /       Appointment p���U  ����U  ��This_stuffs_This_stuffs_ �U  @���U  ����U  ����U   ���U  �VT��  �x /       Some_stuffs  ���U  ����U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ����  �x /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �����  Y�x /       Some_stuffs ����U  ����U   �This_stuffs_This_stuffs_ �U  Ћ��U  ����U   ���U  ����U  �\|��  ��x /      Birthday fs �s��U   t��U  �tSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �x��U  <� ��  �y /      Some_stuffs ���U  ����U  ��justforfun_justforfun_ ��U  ����U  @���U  0���U   ���U  I�(��  � y /       Appointment �W��U  �X��U  @Yjustforfun_justforfun_ ��U  @\��U   ]��U  �]��U  �n��U  �̥��  �@y /       Birthday    ���U  p��U  0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �!��U  ��;��  kgy /       Meeting �U  0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  B.[��  hoy /       Workout     ����U  @���U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0���U  ��[��  �oy /      Meeting                        Some_stuffs_Some_stuffs_                                     �����  D�y /       Some_stuffs p���U  ����U  p�This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  ����U  �����  N�y /       Appointment ���U   ��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  ڀ���  w�y /       Appointment @���U  ����U  ��This_stuffs_This_stuffs_ �U   ���U  ����U  @ ��U   ��U  �4���  (�y /      Workout                        justforfun_justforfun_                                       ّ���  �y /       Some_stuffs  ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  i�r��  �y /       Birthday    ����U  `���U  ��Some_stuffs_Some_stuffs_ �U  ���U  `��U  ��U  ���U  �w��  �y /      Workout     �c��U  �d��U  0eSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pj��U  z���  ��y /       Birthday    г��U  p���U  p�Some_stuffs_Some_stuffs_ �U  ����U  p���U  0���U  ���U  �u���  Ļy /       Some_stuffs `h��U   i��U  �iSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  p�*�  e� /       Some_stuffs ���U  ����U  `�This_stuffs_This_stuffs_ �U  `���U  ���U  ����U  ����U  ��A�  �j� /      Some_stuffs  ��U  ���U  `Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  �<��  ��� /       Birthday    ����U  0���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  e���  ��� /      Meeting     ����U  ���U  ��justforfun_justforfun_ ��U  ����U  ���U  ����U  ���U  I_�  ��� /       Meeting ent @g��U  �g��U  �hThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   m��U  t�m�  ʷ� /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ����  �ۄ /      Appointment ����U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ���  #�� /       Meeting     0E��U  �E��U  pFjustforfun_justforfun_ ��U  �H��U  �I��U  0J��U  �J��U  4���  b� /      Meeting �U  �7��U  `8��U   9This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �=��U  4�%�  b(� /      Meeting     ����U  P���U  ЪSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ys-�  [*� /       Meeting     �		��U  `
	��U  �
	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �	��U  ����  �Q� /       Meeting     p���U  ���U  p�This_stuffs_This_stuffs_ �U  ���U  ����U  p���U  0���U  ����  �S� /      Some_stuffs 0J��U  �J��U  �Kjustforfun_justforfun_ ��U  @^��U  �^��U  �O��U  pP��U  ��`	�  y� /       Appointment ���U  ����U  `�justforfun_justforfun_ ��U  ����U  @���U   ���U  ����U  ��e	�  Pz� /       Workout                        This_stuffs_This_stuffs_                                     @ g	�  �z� /       Some_stuffs                    Some_stuffs_Some_stuffs_                                     �Xl	�  �{� /      Workout �U  0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  ���	�  %�� /       Birthday    �`��U  `a��U   bjustforfun_justforfun_ ��U  `d��U  �d��U  �e��U  `f��U  �-
�  ��� /      Some_stuffs ����U  ����U  `�justforfun_justforfun_ ��U   ���U  ����U  `���U   ���U  j�
�  Q�� /       Some_stuffs ����U  `���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  t��
�  �ƅ /      Birthday    ����U  `���U   �This_stuffs_This_stuffs_ �U  ����U  `���U   ���U  ����U  ri�
�  Fǅ /       Birthday    л��U  ����U  ��This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  p���U  ���
�  ZɅ /       Appointment �U��U  �V��U  P[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �l��U  Dt&�  ,� /      Workout     �6��U   7��U  �7justforfun_justforfun_ ��U  P9��U  �9��U  p:��U  0;��U  I,��  �� /       Workout     �9��U  �:��U  p;justforfun_justforfun_ ��U  �>��U  ?��U  �?��U  P@��U  .ֽ�  �� /      Birthday    ���U  ����U  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ����  �� /       Meeting     �`��U  �a��U  `fjustforfun_justforfun_ ��U  �g��U  �h��U  pj��U  0k��U  TK�  8� /       Some_stuffs 0���U  ����U  p�Some_stuffs_Some_stuffs_ �U  ����U  ����U  p���U  ����U  K�K�  =8� /       Appointment PL��U  M��U  �MThis_stuffs_This_stuffs_ �U  �P��U  Q��U  �Q��U  PR��U  9cQ�  �9� /       Birthday    �<��U  �=��U   >This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �A��U  ͰU�  �:� /       Meeting     P���U  ����U  P�Some_stuffs_Some_stuffs_ �U  ����U  P���U  ����U  ����U  ��W�  N;� /       Meeting     ����U  0��U  ��This_stuffs_This_stuffs_ �U  ����U  p���U  0���U  ����U  ��[�  i<� /      Meeting ffs ���U  ����U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  y{��  [_� /       Workout     @ ��U  � ��U  @!justforfun_justforfun_ ��U  �#��U  �$��U   %��U  �%��U  j���  �`� /       Some_stuffs �L��U  �M��U  @NThis_stuffs_This_stuffs_ �U  �P��U   Q��U  �Q��U   R��U  ���  ub� /       Meeting     ����U  @���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  5��   c� /       Some_stuffs 0e��U  �e��U  �fSome_stuffs_Some_stuffs_ �U  �i��U  pj��U  0k��U  �k��U  a�  Jh� /       Birthday    ���U  ����U   �justforfun_justforfun_ _ �U   ���U  ����U   ���U  ����U  �͗�  C�� /       Meeting      ���U  ����U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  rP�  ��� /       Some_stuffs ����U  @���U  ��justforfun_justforfun_ ��U  0���U  ����U  0���U  ����U  ��  ^�� /      Some_stuffs ���U  ����U  P�Some_stuffs_Some_stuffs_ �U  @���U  ���U  ���U  ����U  ��5�  ��� /       Meeting     �P��U  �Q��U  pRThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   W��U  ���  :Ն /       Workout     Ц��U  ����U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  LG��  �׆ /      Workout     `���U   ���U  ��justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  `���U  �:��  a؆ /       Workout     ����U  p���U  0�This_stuffs_This_stuffs_ �U  ����U  0���U  ����U  ����U  ���  �چ /       Appointment  b��U  �b��U   cSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �g��U  �7��  �چ /       Workout     �;��U  `<��U  �<This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  PO��U  L�L�  !�� /      Meeting     ���U  ����U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  �L��  �"� /       Appointment ����U  P���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  ����  �'� /       Workout �U  �`��U  �a��U  bjustforfun_justforfun_ ��U  �d��U  Pe��U   f��U  �f��U  S��  �)� /      Workout     0���U  ����U  ��Some_stuffs_Some_stuffs_ �U  p���U  0���U  ����U  ����U  z�~�  {K� /       Workout     ����U  ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  W��  `L� /       Appointment 0��U  ���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0��U  �b��  cL� /       Birthday    ����U  0���U  ��Some_stuffs_Some_stuffs_ �U  ����U  p���U  0���U  ����U  䲒�  �P� /      Appointment ��U  ���U  �Some_stuffs_Some_stuffs_ �U  ���U  ���U  p��U  0��U  U��  q� /      Workout     ����U  0���U  P
justforfun_justforfun_ ��U  ����U   ���U  ����U  @���U  (��  �r� /       Meeting �U  ����U  ����U  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P��U  A���  ș� /       Some_stuffs p���U   ���U  ��Some_stuffs_Some_stuffs_ �U  ����U  P���U  ����U  ����U  �:��  >�� /      Birthday     E��U  �F��U  0KThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  \��U  �G�  y�� /      Birthday    p���U  0���U  ��justforfun_justforfun_ ��U  P���U  ���U  ����U  P���U  Q.J�  �� /       Workout ent 0>��U  �>��U  p?Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  �B��U  !���  �� /       Meeting ffs @0��U  �0��U  �1This_stuffs_This_stuffs_ �U  �3��U  p4��U  5��U  �5��U  ����  g� /      Meeting     @^��U  �^��U  �OSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  pT��U  �1u�  �� /      Some_stuffs `���U   ���U  ��Some_stuffs_Some_stuffs_ �U  ����U  `���U   ���U  ����U  [�{�  G� /       Birthday    �n��U  �o��U  @pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �t��U  ��  j� /       Appointment ��U  ���U  �justforfun_justforfun_ _ �U  ���U  ���U  p��U  0��U  �ؕ�  �� /       Appointment @���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  -�  �8� /       Birthday    ����U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  d%�   9� /      Some_stuffs ����U  `���U  `�This_stuffs_This_stuffs_ �U   ���U  ����U  `���U   ���U  ���  �[� /       Workout �U  �j��U  `k��U  �kSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   p��U  ����  �^� /      Meeting      ���U  ����U  `�Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   ���U  �O�  �� /       Workout     ����U  `���U  ��Some_stuffs_Some_stuffs_ �U  ����U  `���U  е��U  ����U  �YT�  H�� /      Meeting     0���U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  M��  �� /      Birthday    ����U  p���U  �justforfun_justforfun_ ��U  ����U  0���U  ����U  p���U  ����  쫈 /       Meeting     ����U  `���U  ��Some_stuffs_Some_stuffs_ �U  ���U  `��U  ��U  ���U  �9��  k�� /       Meeting     ����U  ����U  ��justforfun_justforfun_ ��U  ����U  @���U   ���U  ����U  �l��  x�� /       Meeting     ���U  й��U  P�justforfun_justforfun_ ��U  ����U  P���U  ���U  ����U  �e��  ı� /       Appointment ���U  0 ��U  � Some_stuffs_Some_stuffs_ �U  0$��U  �$��U  �%��U  0&��U  �m��  �؈ /      Meeting                        This_stuffs_This_stuffs_                                     �e�@�  �� /      Appointment ���U  ����U  P�justforfun_justforfun_ ��U  @���U  ���U  ���U  ����U  zgA�  �Г /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             r�tA�  &ԓ /       Appointment `���U   ���U  ��justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  `���U  �-uA�  Eԓ /       Birthday    pm��U  0n��U  �nSome_stuffs_Some_stuffs_ �U  pq��U  �q��U  pr��U  �r��U  i�yA�  qՓ /       Appointment ����U  @���U  �justforfun_justforfun_ ��U  P���U  ���U   ���U  ����U  ���A�  o�� /       Workout     @_��U  P���U  �`Some_stuffs_Some_stuffs_ �U  �b��U  @c��U  �c��U  �d��U  ���A�  E�� /       Appointment ���U  p��U  0Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ���U  EB�  ��� /      Meeting     ���U  p���U  �This_stuffs_This_stuffs_ �U  p���U  ���U  p���U   ���U  (}B�  I�� /       Workout     �<��U  �=��U   >Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �A��U  |P�B�  � /      Appointment  4��U  �4��U  `5This_stuffs_This_stuffs_ �U  �7��U  `8��U   9��U  �9��U  �ʡB�  :!� /       Appointment p��U  ���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ���C�  �j� /      Meeting     @���U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  	��C�  �j� /       Some_stuffs �p��U  �q��U  0rSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0w��U  �1TD�  o�� /      Some_stuffs p���U  ����U  p�justforfun_justforfun_ ��U  � 	��U  @	��U  �	��U  @	��U  (WD�  )�� /       Birthday    @X��U  �X��U  �Yjustforfun_justforfun_ ��U  @\��U  �\��U  @]��U   ^��U   1�D�  ��� /       Meeting ent ��U  ���U  This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  P��U  UQ�D�  ��� /      Appointment ����U   ���U  ��This_stuffs_This_stuffs_ �U  `���U   ���U  ����U  ����U  ��E�  ��� /       Some_stuffs P���U  ���U  ЦSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �x�E�  ��� /       Some_stuffs ���U  ���U   justforfun_justforfun_ ��U  @
��U  �
��U  @��U   ��U  ⇑E�  �� /       Appointment �`��U  `a��U   bThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `f��U  �q�E�  �� /      Some_stuffs ����U  `���U  ��justforfun_justforfun_ _ �U  ����U   ���U  ����U  @���U  �%F�  �� /       Birthday    �Y��U  0Z��U  �ZSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  �^��U  ��4F�  n� /       Workout     л��U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  *�7F�  I� /       Meeting     0���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  p���U  ����U  p���U  )P�F�  ).� /       Meeting     ���U  ���U  0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @��U  ���F�  75� /       Some_stuffs P���U  ���U  иSome_stuffs_Some_stuffs_ �U  ����U  P���U  м��U  P���U  x�YG�  {V� /       Some_stuffs ���U  0��U  �Some_stuffs_Some_stuffs_ �U  p��U  0��U  ���U  0��U  ��H�  E�� /      Meeting      ���U  ����U   �Some_stuffs_Some_stuffs_ �U  `���U  ���U  ����U  ���U  �H�  ��� /       Some_stuffs ���U  ���U  0Some_stuffs_Some_stuffs_ �U  ���U  @��U  ���U  @��U  ��H�  ã� /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             l�5I�  UЕ /      Appointment �*��U  P+��U  �+Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �/��U  ��:I�  �ѕ /       Birthday    �3��U  p4��U  5justforfun_justforfun_ _ �U  �7��U  P8��U  �8��U  �9��U  ��I�  �� /      Some_stuffs �9��U  �:��U  p;This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P@��U  ��I�  �� /       Meeting ffs ����U  P���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ���I�  �� /       Meeting     |��U  �|��U  �}This_stuffs_This_stuffs_ �U  ���U  P���U  ���U  ����U  ��I�  �� /       Appointment p���U  ���U  p�Some_stuffs_Some_stuffs_ �U  ���U  ����U  p���U  0���U  �PYJ�  �� /       Meeting     ���U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  M�jJ�  a� /      Meeting     ����U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  	�-L�  Ւ� /       Some_stuffs ���U  0��U  �Some_stuffs_Some_stuffs_ �U  p��U  0��U  ���U  0��U  �U/L�  I�� /      Appointment  $��U  �%��U   +Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �:��U  (I�L�  ɳ� /       Birthday    д��U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �ڳL�  6�� /       Appointment 0���U  ����U  0�This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  �~OM�  ݖ /       Birthday U  0F��U  �F��U  pGThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  pK��U  a,QM�  |ݖ /       Meeting      ���U  ����U  ��This_stuffs_This_stuffs_ �U  0���U  ����U  ����U  p���U  �=TM�  Eޖ /      Workout  nt P���U  Щ��U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0���U  l
�M�  � /      Appointment  E��U  �F��U  0KThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  \��U  ��M�  � /       Birthday     ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  p���U  ���U  ж��U  ���N�  �+� /      Some_stuffs 0���U  ����U  �justforfun_justforfun_ ��U  p���U  ����U  p���U  0���U  ��O�  XR� /       Appointment  E��U  �F��U  0KThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  \��U  �&O�  �U� /       Appointment ����U  0���U  �Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ���U  ��-O�  rW� /      Workout     ����U  ����U  НSome_stuffs_Some_stuffs_ �U  0���U  ���U  p���U  0���U  ���O�  �~� /       Meeting     `���U   ���U  �justforfun_justforfun_ ��U  ����U  ����U  ����U  @���U  ą�O�  � /      Birthday    Н��U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��HP�  ��� /       Appointment и��U  ����U  P�This_stuffs_This_stuffs_ �U  м��U  P���U  ���U  о��U  ��PP�  �� /       Appointment                    Some_stuffs_Some_stuffs_                                     �SP�  ʢ� /       Meeting     ���U  p���U  0�This_stuffs_This_stuffs_ �U  p���U  ���U  ����U  p���U  �@UP�  #�� /       Some_stuffs ����U  @���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  I��P�  �ŗ /       Birthday    ����U  @���U  �Some_stuffs_Some_stuffs_ �U  P���U  ���U   ���U  ����U  4�P�  �ŗ /      Birthday U  ����U  ����U  p�This_stuffs_This_stuffs_ �U  ����U  @���U  ����U  ����U  :��P�  Ǘ /       Appointment  c��U  �c��U  `dThis_stuffs_This_stuffs_ �U  �f��U  �g��U  `h��U   i��U  ,K�P�  	ɗ /       Birthday    @'��U   (��U  �(Some_stuffs_Some_stuffs_ �U  �+��U   ,��U  �,��U  �-��U  sz�P�  �˗ /       Appointment ���U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  l�R�  5� /      Workout     pF��U  0G��U  �GSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  0L��U  )fR�  �� /       Some_stuffs 0���U  ����U  p�This_stuffs_This_stuffs_ �U  ����U  0���U  ����U  0���U  2R�R�  ><� /       Meeting     �+��U   ,��U  �,This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �1��U  DA�R�  L?� /      Birthday nt �(��U  �)��U  @*Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �.��U  y��R�  ;B� /       Workout �U  �l��U  `m��U   justforfun_justforfun_ ��U  �p��U  �q��U  0r��U  �r��U  ,l|�  �� /      Workout     ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  ����U  P���U  ����U  a�r|�  <� /       Some_stuffs �i��U  pj��U  0kThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  po��U  �}�  �� /       Some_stuffs ����U  P���U  �Some_stuffs_Some_stuffs_ �U  P���U  ����U  ����U  P���U  ��}�  	8� /      Meeting     p ��U  0��U  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0��U  �֘}�  �9� /       Meeting ffs `���U   ���U  ��Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U   ���U  �H�}�  �;� /       Workout     ���U  ����U  `�This_stuffs_This_stuffs_ �U  ����U  `���U  ���U  ����U  0��}�  �>� /       Meeting �U  ����U  @���U  P�justforfun_justforfun_ ��U  P���U  Т��U  ����U  P���U  �,~�  j_� /       Workout     ����U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �C6~�  �a� /      Some_stuffs �z��U  `{��U   |Some_stuffs_Some_stuffs_ �U  p��U  0���U  ����U  ����U  R�C~�  Re� /       Birthday    p���U  ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U   k�~�  4�� /       Some_stuffs ����U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��~�  `�� /       Some_stuffs  V��U  �V��U  �Wjustforfun_justforfun_ ��U  �Y��U  0Z��U  �Z��U  0[��U  ���~�  b�� /       Appointment 0���U  ����U  p�Some_stuffs_Some_stuffs_ �U  ����U  p���U  ����U  p���U  e�~�  ��� /       Appointment `:��U   ;��U  �;Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   @��U  ���~�  :�� /      Meeting     p��U  0��U  0justforfun_justforfun_ ��U   +��U  �+��U  �/��U  p0��U  �8o�  ��� /       Appointment  ���U  ����U  �rThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �w��U  ��v�  볣 /       Meeting      ��U  ���U   Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   #��U  ����  �ң /       Appointment �G��U  0H��U  �HSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  �M��U  vM��  �ӣ /      Birthday    �2��U   3��U   4Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `8��U  ���  �֣ /       Birthday    ���U  й��U  P�This_stuffs_This_stuffs_ �U  ����U  P���U  ���U  ����U  a���  \ۣ /       Birthday    P���U  ����U  P�This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  ����U   C���  4�� /       Some_stuffs ����U  `���U  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  Kݎ��  ��� /       Meeting ffs �F��U   G��U  �GThis_stuffs_This_stuffs_ �U  �I��U  @J��U  �J��U  @K��U  �ꑀ�  e�� /       Meeting     �<��U  0=��U  �=Some_stuffs_Some_stuffs_ �U  p@��U  �@��U  pA��U  �A��U  hw���  ` � /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             i����  �� /       Workout      c��U  �c��U  `dThis_stuffs_This_stuffs_ �U  �f��U  �g��U  `h��U   i��U  I�0��  %� /       Meeting     ����U  `���U  ��justforfun_justforfun_ ��U  ���U  `��U  ��U  ���U  �}7��  �&� /      Appointment p���U  0���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �>��  �(� /       Some_stuffs                    justforfun_justforfun_                                       1�Ɂ�  >L� /       Some_stuffs 0f��U  �g��U  �ijustforfun_justforfun_ ��U  �p��U  �q��U  �s��U  �t��U  Dn΁�  lM� /      Meeting     `���U  ����U  `�This_stuffs_This_stuffs_ �U  ����U   ���U  ����U  `���U  :�ρ�  �M� /       Some_stuffs ����U  @���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��R��  Qo� /      Workout     е��U  ����U  �Some_stuffs_Some_stuffs_ �U  ����U  ����U  ���U  ����U  	%]��  �q� /       Birthday    ����U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  p��  ��� /       Some_stuffs ����U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  }����  ߽� /      Birthday    ���U  ����U  0�This_stuffs_This_stuffs_ �U   ���U  ����U  ����U  @���U  �酃�   /       Workout      o��U  �o��U  �pThis_stuffs_This_stuffs_ �U  Ps��U  t��U  �t��U  �u��U  2u���  �� /       Some_stuffs 0���U  ����U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  3!���  �ä /       Some_stuffs                    justforfun_justforfun_ _Some_stuffs_Some_stuffs_             �"��  � /       Workout     ����U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ��4��  �� /      Appointment P��U  ���U  PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p#��U  Ђ5��  �� /       Appointment ���U  ����U  0�Some_stuffs_Some_stuffs_ �U   ���U  ����U  ����U  @���U   nɄ�  �� /       Birthday    ���U  ����U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  ��ʄ�  $� /       Some_stuffs @_��U  P���U  �`This_stuffs_This_stuffs_ �U  �b��U  @c��U  �c��U  �d��U  kτ�  1� /       Some_stuffs ���U  @���U  �justforfun_justforfun_ ��U  @���U  ���U  p���U  ���U  mф�  �� /      Workout �U  0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  40҄�  �� /       Workout     `���U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  �Dc��  "8� /       Birthday    �g��U  �h��U  pjThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �o��U  
�c��  58� /       Workout     ���U  ����U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  �l��  �:� /      Birthday    �O��U  pP��U  �PSome_stuffs_Some_stuffs_ �U  �S��U  pT��U  0U��U  �U��U  ����  �\� /      Birthday U  ��U  ���U  PSome_stuffs_Some_stuffs_ �U  ���U  P��U  ���U  �	��U  kq���  q�� /       Some_stuffs ����U  `���U   �Some_stuffs_Some_stuffs_ �U  ����U  p���U  0���U  ����U  ^Ō��  K�� /      Meeting     ����U  `���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `���U  p���  f�� /       Appointment 0���U   ���U  @�This_stuffs_This_stuffs_ �U  p���U  0���U  ����U  `���U  �蕆�  ��� /       Some_stuffs л��U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  �l&��  ��� /       Workout     0e��U  �e��U  �fThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �k��U  ����  �Υ /      Some_stuffs  ���U  ����U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  x0���  {ҥ /       Meeting     ���U  0��U  �This_stuffs_This_stuffs_ �U  ���U  ���U  p��U  0��U  b!S��  ��� /       Some_stuffs �Q��U  PR��U  �RSome_stuffs_Some_stuffs_ �U  PU��U  �U��U  �q��U  `r��U  ��T��  �� /       Birthday nt  ��U  ���U  0This_stuffs_This_stuffs_ �U   ��U  ���U   ��U  ���U  t�Z��  ��� /      Birthday                       Some_stuffs_Some_stuffs_                                     X���  �!� /       Some_stuffs P[��U  \��U  �`Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �h��U  �v���  �$� /       Workout      ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  �2w��  aC� /       Meeting     p��U  0��U  �justforfun_justforfun_ _ �U  p��U  0��U   &��U  �&��U  Rِ��  �I� /       Meeting     ����U  @���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  5���  �J� /      Meeting     p ��U  0��U  pSome_stuffs_Some_stuffs_ �U  0��U  ���U  p��U  0��U  ���  �m� /      Meeting     ����U  P���U  �Some_stuffs_Some_stuffs_ �U  ����U  ����U  0���U  ����U  MN���  A�� /      Birthday U  PL	��U  M	��U  �M	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Q	��U  �վ��  A�� /       Meeting ent p7��U  08��U  �8Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  >��U  t����  j� /      Meeting     ����U  P���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��z��  �� /      Meeting     @^��U  �^��U  �OSome_stuffs_Some_stuffs_ �U  pR��U  �R��U  �S��U  pT��U  �p���  �� /       Some_stuffs ^��U  �^��U  @_justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  @c��U  yr��  �/� /       Birthday fs P	��U  �	��U  P	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @	��U  �j!��  �3� /      Workout     �{��U  0|��U  �|This_stuffs_This_stuffs_ �U  `���U  ����U  `���U   ���U  |DÍ�  �\� /      Workout ffs @Y��U   Z��U  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   `��U  �����  �*� /       Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �O���  X+� /       Some_stuffs ����U  0���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ����  W� /       Workout �U  ����U  ����U  ��justforfun_justforfun_ ��U  0���U   ���U  @���U   ���U  �����  �X� /      Birthday    p��U  0��U  0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p0��U  ��-��  Nz� /       Meeting     `6��U   7��U  �7Some_stuffs_Some_stuffs_ �U  `:��U   ;��U  �;��U  `<��U  ��7��  �|� /      Some_stuffs �4��U  p5��U  �9justforfun_justforfun_ ��U   E��U  �F��U  0K��U  �K��U  �'>��  �~� /       Some_stuffs 0���U  ����U  p�Some_stuffs_Some_stuffs_ �U  ����U  p���U  ����U  p���U  �HA��  N� /       Some_stuffs �h��U   i��U  �iSome_stuffs_Some_stuffs_ �U  �l��U   m��U  �m��U  @n��U  ��չ�  P�� /      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �F۹�  ��� /       Some_stuffs p��U  ���U  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p��U  <#\��  �ǲ /      Some_stuffs ���U  ����U  ��justforfun_justforfun_ ��U  ����U  @���U  0���U   ���U  	���  �� /       Birthday U  0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  �0���  �� /       Some_stuffs  ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  p���U  P���U  ���U  �����  � /      Meeting     �g��U  �h��U  pjThis_stuffs_This_stuffs_ �U  �m��U  @n��U   o��U  �o��U  {
��  ;�� /       Birthday nt ����U  `���U   �Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  Û��  �� /       Meeting  fs � ��U  �!��U  p"This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   (��U  |Ǩ��  �� /      Appointment                    This_stuffs_This_stuffs_                                     C0���  �d� /       Workout     �R	��U  S	��U  �S	justforfun_justforfun_ 	��U  �U	��U  @V	��U  �V	��U  @W	��U  �rμ�  h� /       Birthday    ����U  @���U  0�Some_stuffs_Some_stuffs_ �U  P���U  ���U  p���U  0���U  UҼ�  �h� /      Some_stuffs 0��U  ���U  �justforfun_justforfun_ ��U  p��U  ���U  ���U  0 ��U  ��ܼ�  �k� /       Some_stuffs 0p��U  �p��U  pqThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Pu��U  �8c��  #�� /       Workout     0���U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  �1j��  쏳 /       Birthday    � 	��U  @	��U  �	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �	��U  ��k��  Y�� /       Some_stuffs                    This_stuffs_This_stuffs_                                     Hg���  ݵ� /       Appointment P[��U  \��U  �`This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �h��U  ����  ��� /      Meeting     ���U   ��U  �justforfun_justforfun_ ��U  p��U  ���U  ���U  @��U  T����  2س /       Appointment 0���U  ����U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  DN���  lٳ /      Some_stuffs �/��U  p0��U  �4This_stuffs_This_stuffs_ �U  �>��U  �?��U   E��U  �F��U  ����  �۳ /       Birthday    ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  �����  �ܳ /       Workout ffs ����U  ����U  `�This_stuffs_This_stuffs_ �U   ���U  ���U  ����U  ���U  N����  �ݳ /       Appointment �0��U  �1��U   2This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �5��U  ���  ޳ /       Birthday U   ��U  ���U   This_stuffs_This_stuffs_ �U   ��U  ���U  `��U  ���U  �J���  �߳ /       Birthday    ���U  ж��U  P�justforfun_justforfun_ ��U  P���U  ���U  ����U  P���U  P+��  �� /       Meeting     ����U   ���U  ��Some_stuffs_Some_stuffs_ �U  е��U  ����U  ���U  й��U  �J+��  �� /       Birthday U  PH��U  I��U  �IThis_stuffs_This_stuffs_ �U  PL��U  M��U  �M��U  �N��U  b0��  � /       Some_stuffs P���U  Ј��U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  �yƿ�  �*� /      Appointment @\��U  �\��U  @]Some_stuffs_Some_stuffs_ �U  �_��U  �`��U   a��U  �a��U  #�ƿ�  �*� /       Meeting     ����U  P���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  ӿ�  �-� /       Appointment `f��U   g��U   lThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �r��U  ��տ�  �.� /       Birthday    `���U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  =Q��  $N� /      Appointment                    justforfun_justforfun_                                       �D\��  �P� /       Birthday    0E��U  �E��U  pFThis_stuffs_This_stuffs_ �U  �H��U  �I��U  0J��U  �J��U  �]��  VQ� /       Meeting     p���U  ����U  ��justforfun_justforfun_ ��U   ���U  ����U  @���U  ����U  ����  �t� /       Workout     `6��U   7��U  �7justforfun_justforfun_ ��U  `:��U   ;��U  �;��U  `<��U  &����  �w� /      Some_stuffs P
��U  �
��U  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  `����  �z� /       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_              ����  ��� /       Meeting �U  �K��U  0L��U  �LSome_stuffs_Some_stuffs_ �U  �O��U  pP��U  �P��U  �Q��U  �:���  ��� /       Some_stuffs �s��U   t��U  �tjustforfun_justforfun_ ��U  w��U  �w��U  x��U  �x��U  �{���  ��� /      Meeting �U  Ъ��U  ����U  P�Some_stuffs_Some_stuffs_ �U  Ю��U  ����U  ���U  ����U  ��"��  CŴ /       Some_stuffs                    Some_stuffs_Some_stuffs_                                     ��*��  aǴ /       Birthday    ����U  ����U  @�Some_stuffs_Some_stuffs_ �U   ���U  ����U  0���U  ����U  p],��  �Ǵ /       Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             v:��  J˴ /      Some_stuffs л��U  ����U  ��This_stuffs_This_stuffs_ �U  0���U  ���U  ����U  p���U  `����  �� /       Some_stuffs ����U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  a����  �� /       Some_stuffs  ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  `���U  ����U  `���U  �����  g� /      Some_stuffs ����U  P���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �_���  �� /       Meeting      &��U  �&��U  0Some_stuffs_Some_stuffs_ �U  0��U  ���U  p��U  ���U  mT��  u� /      Appointment pv��U  0w��U  �wSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0|��U  ��^��  8� /       Meeting     ����U  ���U  ЮSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ����  �7� /      Meeting     P���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �C���  0e� /       Meeting     ����U  p���U  0�justforfun_justforfun_ ��U  ���U  ����U  ����U  @���U  d:��  @�� /      Appointment pF��U  0G��U  �GThis_stuffs_This_stuffs_ �U  0J��U  �J��U  �K��U  0L��U  �((��  N�� /       Workout     �w��U  �x��U  PsThis_stuffs_This_stuffs_ �U  v��U  �v��U  0~��U  �~��U  �,5��  ��� /       Appointment ����U  P���U  ��justforfun_justforfun_ _ �U  ���U  ����U  P���U  ����U  I����  }�� /       Birthday                       This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_             �����  1�� /      Some_stuffs 0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  "����  ��� /       Some_stuffs е��U  ����U  �Some_stuffs_Some_stuffs_ �U  ����U  ����U  ���U  ����U  �#F��  �Ե /       Birthday    ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  �!a��  m۵ /       Birthday nt ����U  @���U  ��Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ���U  m�b��  �۵ /      Meeting �U  г��U  p���U  p�Some_stuffs_Some_stuffs_ �U  ����U  p���U  0���U  ���U  �����  F� /      Birthday nt �2��U  @3��U  �3Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P8��U  @Zx��  �"� /       Birthday U  �H��U  @I��U  �IThis_stuffs_This_stuffs_ �U  �K��U  @L��U  �L��U  �M��U  �az��  m#� /       Meeting     ����U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  �;���  �%� /      Appointment P�	��U  Њ	��U  P�	Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   �	��U  Ѿ���  b(� /       Appointment @���U  ����U  @�This_stuffs_This_stuffs_ �U  ����U  P���U  д��U  P���U  ����  �*� /       Meeting ffs �g��U  �h��U  pjSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �o��U  �G��  \L� /      Workout     ����U  p���U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U   ?���  �p� /       Some_stuffs P[��U  \��U  �`This_stuffs_This_stuffs_ �U   l��U  �l��U  �g��U  �h��U  �ͩ��  q� /      Appointment @��U  ���U  @This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ��U  �Ѵ��  �s� /       Appointment �O��U  pP��U  �Pjustforfun_justforfun_ ��U  �S��U  pT��U  0U��U  �U��U  ��A��  �� /       Birthday fs ����U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  HG��  ]�� /       Meeting ent �t��U  �u��U  vThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `{��U  >V��  ?�� /       Appointment                    This_stuffs_This_stuffs_                                     T�W��  ��� /       Meeting     ���U  @��U  �This_stuffs_This_stuffs_ �U   ��U  ���U  @ ��U  � ��U  ]+a��  �� /      Birthday     ���U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ^���  ��� /       Some_stuffs                    Some_stuffs_Some_stuffs_                                     �����  �¶ /       Birthday    P���U  ���U  ��This_stuffs_This_stuffs_ �U  ���U  ����U  P���U  ���U  1����  ^ƶ /       Birthday nt �z��U  `{��U   |Some_stuffs_Some_stuffs_ �U  p��U  0���U  ����U  ����U  ͌�p,�  Q2 &/      Some_stuffs p���U  ���U  ��justforfun_justforfun_ ��U  ���U  ����U  @���U  ����U  Zp�p,�  '7 &/       Birthday    ����U  ���U  ��justforfun_justforfun_ ��U  ����U  0���U  ����U  `���U  (��p,�  �7 &/       Meeting     ����U  p���U  0�Some_stuffs_Some_stuffs_ �U  ���U  ����U  ����U  @���U  ��iq,�  �\ &/      Workout     @���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��tq,�  d_ &/       Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             -vq,�  �_ &/       Some_stuffs ���U  p���U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  �׀q,�  �b &/       Some_stuffs �(��U  �)��U  @*This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �.��U  ���q,�  �� &/       Birthday nt @t��U  �t��U  �ujustforfun_justforfun_ _This_stuffs_This_stuffs_ �U  Pz��U  ��r,�  � &/       Birthday nt �w��U  px��U  0yjustforfun_justforfun_ _This_stuffs_This_stuffs_ �U  �}��U  Yץr,�  �� &/       Some_stuffs �L��U  �M��U  @^Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  �R��U  ��r,�  � &/      Birthday    ���U  ����U  `�This_stuffs_This_stuffs_ �U  ����U  @���U   ���U  ����U  �Ьr,�  P� &/       Birthday    ����U  P���U  ��This_stuffs_This_stuffs_ �U  ����U  @���U  ����U  ����U  �z+s,�  �� &/      Some_stuffs @	��U  �	��U  �	This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  `	��U  �Ds,�  � &/       Meeting     P���U  ���U  ЦSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ���s,�  I� &/      Workout �U  �	��U    	��U  � 	This_stuffs_This_stuffs_ �U  �"	��U  0#	��U  �#	��U  0$	��U  q�s,�  &� &/       Workout     ���U  ж��U  P�This_stuffs_This_stuffs_ �U  P���U  ���U  ����U  P���U  Tsut,�  6$&/      Meeting ent  ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ж��U  D!u,�  LK&/      Birthday     &��U  �&��U  0This_stuffs_This_stuffs_ �U  0��U  ���U  p��U  ���U  �	�u,�  �k&/      Workout     @(��U  �(��U  p)Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �-��U  *z�u,�  il&/       Birthday    p���U  0���U  ��This_stuffs_This_stuffs_ �U  ���U  ����U  ���U  ����U  �M�u,�  �n&/       Some_stuffs                    justforfun_justforfun_                                       9��u,�  Sr&/       Workout �U  p?��U  �?��U  p@This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �D��U  �=6v,�  �&/       Meeting     p��U  0��U  �Some_stuffs_Some_stuffs_ �U  �	��U  0
��U  �
��U  ���U   <v,�  ��&/       Birthday    е��U  ����U  �Some_stuffs_Some_stuffs_ �U  ����U  ����U  ���U  ����U  2�=v,�  ��&/       Workout ffs  ���U  ����U  ��This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  p���U  ��v,�  +�&/       Birthday    ���U  p���U  0�justforfun_justforfun_ _ �U  ����U  p���U  ����U  p���U  <l�v,�  W�&/      Workout �U  0f��U  �g��U  �iSome_stuffs_Some_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  ���v,�  x�&/       Appointment 0e��U  �e��U  �fSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �k��U  �Mdw,�  n�&/       Meeting                        This_stuffs_This_stuffs_                                     �N�w,�  �	&/       Some_stuffs �8��U  �9��U   :Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �=��U  |��w,�  _
&/      Meeting �U  0f��U  �g��U  �iThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �t��U  q��w,�  f&/       Appointment pv��U  0w��U  �wSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0|��U  䲍x,�  �0&/      Workout                        This_stuffs_This_stuffs_                                     ��!y,�  �V&/       Appointment ����U  � ��U  @This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U   ��U  �y8y,�  H\&/      Meeting                        This_stuffs_This_stuffs_                                     X½y,�  g~&/       Birthday                       justforfun_justforfun_                                       2i�y,�  ��&/       Appointment ����U   ���U  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  UU�y,�  v�&/      Appointment `���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `���U  1�Xz,�  �&/       Meeting     � 	��U  @	��U  �	justforfun_justforfun_ 	��U  �	��U  �	��U  @	��U  �	��U  ��]z,�  c�&/       Some_stuffs ����U  @���U  ��This_stuffs_This_stuffs_ �U   ���U  ����U  @ ��U  � ��U  ���z,�  3�&/      Birthday    @*��U   +��U  �+Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @0��U  H��{,�  }�&/       Meeting     `���U   ���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  *B|,�  i&/       Some_stuffs ����U   ���U  ��This_stuffs_This_stuffs_ �U  @ ��U   ��U  ���U  P��U  )�|,�  �&/       Appointment P���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  P���U  ���U  ����U  <�0|,�  �&/      Meeting �U  0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  *#�|,�  	@&/       Workout     @���U    ��U  �justforfun_justforfun_ ��U  ���U  P��U   ��U  ���U  d=�|,�  B&/       Meeting     е��U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��|,�  �F&/      Meeting     ���U  ����U  P�Some_stuffs_Some_stuffs_ �U  ���U  ����U  ����U  P���U  S�|,�  2G&/       Workout     ����U  0��U  ��This_stuffs_This_stuffs_ �U  ����U  p���U  0���U  ����U  �*�|,�  6G&/       Workout     0���U  ����U  ��This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  !�I},�  �f&/       Meeting                        Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_             �R},�  �h&/      Appointment p��U  0��U  0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p0��U  KQ^},�  l&/       Birthday nt ����U  ����U  p This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  ��_},�  �l&/       Birthday nt  ^	��U  �^	��U   _	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �b	��U  `��~,�  |�&/       Appointment �7��U   8��U  �_justforfun_justforfun_ ��U  p:��U  0;��U  �;��U  0<��U  l/,�  5�&/      Birthday fs 0r��U  �r��U  �sThis_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  px��U  ���,�  �&/      Workout      ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  `���U   ���U  ����U  ��,�  �&/       Some_stuffs  ���U  ����U  ��This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  `���U  Ӊ�,�  B&/       Workout     �0��U  �1��U   2justforfun_justforfun_ _ �U   4��U  �4��U   5��U  �5��U  �ּ,�  b&/       Meeting     `V��U   W��U  �WSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ]��U  `0�,�  �&/       Birthday    P[��U  \��U  �`This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �h��U  ��Y�,�  �/&/      Appointment ����U  P���U  �This_stuffs_This_stuffs_ �U  `���U   ���U  ���U  ����U  мg�,�  "3&/       Birthday     E��U  �F��U  0KSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  \��U  q��,�  fS&/       Workout     `���U   ���U  ��justforfun_justforfun_ ��U  `���U   ���U  ����U  `���U  �G��,�  ^W&/      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ��$�,�  �&/      Workout     ����U  `���U  ��Some_stuffs_Some_stuffs_ �U  ����U  `���U  е��U  ����U  ���,�  .�&/       Birthday    ����U  P���U  �This_stuffs_This_stuffs_ �U  `���U   ���U  ���U  ����U  􉯂,�  ��&/       Workout     ���U  й��U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �ᰂ,�  ��&/       Birthday fs p@��U  �@��U  pAThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �E��U  4��,�  �&/      Birthday U  ��U  ���U  �justforfun_justforfun_ ��U  ���U  ���U  p��U  0��U  ꨱ�,�  !�&/       Some_stuffs p���U  0���U  ��This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  %���,�  ��&/       Some_stuffs @���U  ����U  @�justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  ����U  ��g�,�  �v&/      Appointment �s��U  pt��U  0ujustforfun_justforfun_ ��U  �w��U  px��U  0y��U  �y��U  ��~�,�  �|&/       Workout �U  p���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �g�,�  V�&/       Meeting     л��U  ����U  ��justforfun_justforfun_ ��U  0���U  ���U  ����U  p���U  e�,�  ��&/      Birthday    ����U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  YP�,�  '�&/       Appointment �#��U  p$��U  0%This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   +��U  K��,�  ��&/      Appointment ����U  ����U  p�justforfun_justforfun_ ��U  0���U  ����U  ���U  ����U  ���,�  ,�&/       Some_stuffs ����U  ����U  ��justforfun_justforfun_ _ �U  ����U  @���U   ���U  ����U  �秭,�  ��&/       Some_stuffs ����U  ����U   �justforfun_justforfun_ _ �U  ���U  P��U  ��U  ���U  Ji��,�  �&/       Workout     �P��U   Q��U  �QThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  `U��U  |/9�,�  ��&/      Meeting ffs �O��U  pP��U  �PThis_stuffs_This_stuffs_ �U  �S��U  pT��U  0U��U  �U��U  ,AѮ,�  �&/      Birthday     E��U  �F��U  0Kjustforfun_justforfun_ ��U  �U��U  �V��U  P[��U  \��U  	`Ѯ,�  �&/       Appointment `���U   ���U  ��justforfun_justforfun_ ��U  ����U  @���U   ���U  ����U  �b�,�  �9&/       Birthday     %��U  �%��U  @&Some_stuffs_Some_stuffs_ �U  @(��U  �(��U  p)��U  *��U  �e�,�  �:&/       Appointment PO��U  �O��U  �PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �T��U  99h�,�  s;&/       Birthday                       Some_stuffs_Some_stuffs_                                     D m�,�  �<&/      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             
���,�  u_&/       Some_stuffs ����U   ���U  ��This_stuffs_This_stuffs_ �U   ���U  ����U  ����U   ���U  ���,�  �d&/       Some_stuffs ����U  p���U  0�This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  p���U  <e
�,�  �d&/      Appointment л��U  ����U  ��Some_stuffs_Some_stuffs_ �U  0���U  ���U  ����U  p���U  1z�,�  >e&/       Workout     `���U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  �G��,�  ��&/       Appointment  t��U  �t��U   uSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �x��U  @��,�  ��&/       Some_stuffs ����U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ����,�  ��&/       Birthday    `���U   ���U  ��Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   ���U  ={��,�  ��&/      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �`$�,�  '�&/      Appointment                    Some_stuffs_Some_stuffs_                                     j�0�,�  Q�&/       Meeting     �M��U  �N��U  POjustforfun_justforfun_ ��U  �Q��U  PR��U  �R��U  PS��U  �o5�,�  ��&/       Birthday     E��U  �F��U  0KSome_stuffs_Some_stuffs_ �U  �U��U  �V��U  P[��U  \��U  �T��,�  O�&/       Meeting     �,��U  �-��U  @.Some_stuffs_Some_stuffs_ �U   1��U  �1��U  �2��U   3��U  �jǱ,�  ��&/       Birthday    ����U  ����U  p This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  � Ա,�  %�&/       Appointment ����U  ����U  `�Some_stuffs_Some_stuffs_ �U   ���U  ����U  `���U   ���U  ��a�,�  k�&/       Birthday    �{	��U  �|	��U  @}	Some_stuffs_Some_stuffs_ �U  �	��U   �	��U  ��	��U   �	��U   �t�,�  4&/       Some_stuffs @b��U  �b��U  �cjustforfun_justforfun_ _ �U  @f��U  �f��U  @g��U  �g��U  ��,�  �(&/      Birthday     ���U  ����U  �rThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �w��U  *K�,�  	)&/       Workout     ����U  ���U  ЮThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  �r�,�  a+&/       Some_stuffs                    justforfun_justforfun_                                       J3��,�  ]M&/       Meeting     @��U   ��U  �This_stuffs_This_stuffs_ �U  ���U  @��U   ��U  ���U  Xї�,�  �M&/       Meeting ffs 0f��U  �g��U  �ijustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  �t��U  U蝳,�  VO&/      Birthday    �e��U  `f��U  �fThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   l��U  �p*�,�  Ps&/       Workout     ����U  ���U  ��justforfun_justforfun_ ��U  ����U  @���U  ����U  @���U  H+>�,�  ]x&/       Workout     p?��U  �?��U  p@This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �D��U  4Է�,�  ��&/      Appointment 0���U   ���U  @�Some_stuffs_Some_stuffs_ �U  p���U  0���U  ����U  `���U  yXǴ,�  {�&/       Birthday fs  ���U  ����U  ��This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  p���U  "1ɴ,�  ��&/       Birthday    @���U  ����U  `�Some_stuffs_Some_stuffs_ �U  ����U  `���U  ����U  `���U  �UV�,�  �&/       Appointment �K��U  @L��U  �Ljustforfun_justforfun_ _ �U  pO��U  �O��U  �P��U   Q��U  �}_�,�  n�&/       Workout     �=��U  �>��U  p?Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pC��U  d�h�,�  ��&/      Workout ent �s��U  pt��U  0uSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  �y��U  ʢm�,�  �&/       Workout ffs  ��U  ���U  @ Some_stuffs_Some_stuffs_ �U  @"��U   #��U  �#��U  �$��U  �	�,�  ��&/       Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ���,�  e�&/       Workout     @���U   ���U  ��Some_stuffs_Some_stuffs_ �U  ����U  @���U   ���U  ����U  6*��,�  B�&/      Birthday    ����U  P���U  ��justforfun_justforfun_ ��U  P���U  ����U  P���U  ����U  +߄�,�  �&/       Appointment ����U  `���U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ���,�  &/      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ғ��,�  �&/       Workout     Ю��U  ����U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  iE��,�  �&/       Appointment p��U  0��U  0Some_stuffs_Some_stuffs_ �U   +��U  �+��U  �/��U  p0��U  �%�,�  �6&/      Workout  U  �	��U  @	��U  �	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �	��U  ��,�  �\&/      Birthday    0���U  ����U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  �r��,�  �]&/       Some_stuffs ����U  `���U  ��This_stuffs_This_stuffs_ �U  ���U  `��U  ��U  ���U  qǷ,�  `&/       Birthday    ���U   ��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @��U  ��O�,�  �&/       Meeting     ����U  0���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  JS�,�  �&/       Some_stuffs `���U  ����U  `�This_stuffs_This_stuffs_ �U  `���U   ���U  ����U   ���U  4~Z�,�  &/      Some_stuffs ���U  P��U   Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  QDn�,�  Ҋ&/       Workout      ��U  ���U  `oSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pt��U  ����,�  ~�&/      Some_stuffs ���U  0 ��U  � Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  0&��U  �惹,�  ��&/      Some_stuffs �	��U  �
��U   justforfun_justforfun_ ��U  @��U  ���U  @��U  ���U  ���,�  �&/       Workout     ����U  @���U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U   &��,�  �&/       Workout �U  0K��U  �K��U  �PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �a��U  �	��,�  �&/       Birthday    ���U  ����U  �justforfun_justforfun_ ��U  ����U  ���U  Ѕ��U  ����U  �!�,�  Y�&/      Workout     ����U  `���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  q7�,�  ��&/       Workout     ����U  ����U  �justforfun_justforfun_ ��U  ����U  `���U  @���U  ���U  �Y��,�  � &/      Birthday    w��U  �w��U  xSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �|��U  h;˺,�  �%&/       Appointment  ���U  ����U  ��justforfun_justforfun_ ��U  ����U  `���U   ���U  ����U  X�O�,�  �G&/       Appointment @\��U  �\��U  @]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �a��U  Х�,�  �n&/       Birthday U   9��U  �9��U  `:This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �>��U  Y�,�  �o&/       Appointment 0~��U  ����U  `�Some_stuffs_Some_stuffs_ �U  ����U  `���U   ���U  ����U  ����,�  o�&/       Meeting ffs �Z��U  0[��U  �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  Lֆ�,�  A�&/      Appointment 0f��U  �g��U  �ijustforfun_justforfun_ ��U  �p��U  �q��U  �s��U  �t��U  �U��,�  �&/       Birthday    0F��U  �F��U  pGSome_stuffs_Some_stuffs_ �U  �I��U  pJ��U  �J��U  pK��U  
��,�  �&/       Appointment ����U   ���U  ��Some_stuffs_Some_stuffs_ �U  ����U  p���U  ����U  p���U  ሚ�,�  L�&/       Birthday    0���U   ���U  @�This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  `���U  ���,�  g�&/      Meeting     ����U  `���U  ��Some_stuffs_Some_stuffs_ �U  ����U  `���U  е��U  ����U  ���,�  d�&/      Appointment �c��U  @d��U  �dSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   i��U  ɖ��,�  ��&/       Workout     0��U  ���U  �Some_stuffs_Some_stuffs_ �U  0"��U  �<��U  0$��U  �$��U  �5�,�  n&/       Appointment ���U  Ш��U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ʿ?�,�  -
&/       Meeting �U  ���U  @��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �E��U  � F�,�  �&/      Birthday nt ����U  P���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ���,�  �/&/      Appointment p��U  0��U   &Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ��b�,�  �T&/       Workout                        justforfun_justforfun_                                       !Vd�,�  U&/       Appointment ����U  p���U  0�Some_stuffs_Some_stuffs_ �U  ����U  0���U  ���U  ����U  ~!t�,�  Y&/      Workout  U  p���U  0���U  ��justforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U  ���U  b��,�  �{&/       Meeting     p���U  0���U  ��Some_stuffs_Some_stuffs_ �U  p���U  ����U  ����U  0���U  ��,�  ��&/      Meeting     0���U  ����U  p�This_stuffs_This_stuffs_ �U  ���U  ����U  P���U  ���U  ��,�  ?�&/       Appointment ���U  @��U   This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �!��U  m9��,�  u�&/      Meeting     @g��U  �g��U  �hThis_stuffs_This_stuffs_ �U   k��U  �k��U  �l��U   m��U  躩�,�  a�&/       Some_stuffs �|��U  �}��U  0~justforfun_justforfun_ ��U  `���U   ���U  ����U  `���U  IE7�,�  ��&/       Workout     @	��U  �@	��U  A	justforfun_justforfun_ 	��U  PC	��U  �C	��U  �D	��U  E	��U  <�F�,�  ��&/      Birthday    @.��U  �.��U  �/Some_stuffs_Some_stuffs_ �U  �2��U   3��U   4��U  �4��U  $���,�  ��&/      Some_stuffs p��U  0��U  0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p0��U  ���,�  ��&/       Appointment Р��U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ���,�  N�&/       Some_stuffs  >��U  �>��U  `?Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pC��U  ��Y�,�  � &/      Some_stuffs  f��U  �f��U   gThis_stuffs_This_stuffs_ �U   i��U  �i��U  �j��U  `k��U  �,b�,�  " &/       Meeting     `���U   ���U  ��Some_stuffs_Some_stuffs_ �U  `���U   ���U  ����U  `���U  2��,�  �> &/       Birthday     �	��U  ��	��U  0�	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �	��U  �z��,�  a@ &/       Birthday    `���U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  ��,�  �C &/      Appointment �P��U  �Q��U  pRSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   W��U  ���,�  j &/       Birthday    ����U  p���U  0�Some_stuffs_Some_stuffs_ �U  ����U  0���U  ����U  ����U  �Ϟ�,�  1j &/      Appointment @��U   ��U  �This_stuffs_This_stuffs_ �U  @��U   ��U  ���U   ��U  �&�,�  Ќ &/       Meeting �U  p ��U  0��U  pThis_stuffs_This_stuffs_ �U  0��U  ���U  p��U  0��U  }F;�,�  ?� &/      Workout     �2��U   3��U   4Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `8��U  !h��,�  T� &/       Some_stuffs 00��U  �0��U  p1justforfun_justforfun_ ��U  04��U  �4��U  05��U  �5��U  kJ��,�  � &/       Appointment �5	��U   6	��U  �6	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `:	��U  "U��,�  t� &/       Appointment `���U   ���U  ��Some_stuffs_Some_stuffs_ �U  `���U  ����U  `���U   ���U  D���,�  ̻ &/      Birthday    p��U  0��U  �Some_stuffs_Some_stuffs_ �U  ���U  ���U  p��U  ���U  ��c�,�  /� &/       Birthday fs `���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��p�,�  �� &/       Workout     Н��U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ,�s�,�  M� &/      Birthday U   ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ����,�  � !&/       Birthday    @���U   ���U  ��This_stuffs_This_stuffs_ �U  ����U  @���U   ���U  p���U  ���,�  a!&/       Meeting                        Some_stuffs_Some_stuffs_                                     ����,�  !&/      Meeting                        Some_stuffs_Some_stuffs_                                     Z��,�  '!&/       Birthday U  �w��U  px��U  0ySome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  �}��U  !���,�  �(!&/       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             R���,�  �*!&/       Birthday    ����U  ���U  ��justforfun_justforfun_ ��U  ����U  0���U  ����U  0���U  x[��,�  [+!&/       Birthday    ����U  `���U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �
-�,�  6S!&/       Birthday     W��U  �W��U  @XThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �\��U  �x��,�  )w!&/      Birthday    ��U  ���U  �justforfun_justforfun_ ��U  ���U  ���U  p��U  0��U  4�M�,�  "�!&/      Appointment                    This_stuffs_This_stuffs_                                     Dc��,�  ��!&/      Birthday                       This_stuffs_This_stuffs_                                     ���,�  7�!&/       Workout     ����U  0��U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ���,�  �"&/       Birthday    ����U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  �.��,�  d9"&/       Meeting     ����U  P���U   �justforfun_justforfun_ ��U  @��U  ���U  ����U  0���U  ����,�  (?"&/      Some_stuffs  E��U  �F��U  0KThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  \��U  �q��,�  �?"&/       Birthday    ����U  p���U  �justforfun_justforfun_ ��U  ���U  й��U  P���U  ���U  ���,�  �?"&/       Appointment `���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �K�,�  @a"&/       Birthday    �;��U  `<��U  �<This_stuffs_This_stuffs_ �U  `?��U   @��U  �N��U  PO��U  �L�,�  �a"&/       Birthday    ����U  p���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  �Gj�,�  i"&/      Meeting      ���U  ����U  ��justforfun_justforfun_ ��U  Н��U  ����U  ����U  p���U  W��,�  �"&/      Birthday    ����U  P���U  �Some_stuffs_Some_stuffs_ �U  ���U  ����U  ����U  ����U  � �,�  ��"&/       Meeting                        This_stuffs_This_stuffs_                                     ���,�  {�"&/      Some_stuffs P���U  ����U  @This_stuffs_This_stuffs_ �U  ����U  ����U  p���U  ����U  �� �,�  9�"&/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             y�$�,�  [�"&/       Birthday    ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  ����U  ����U  ����U  �$&�,�  ��"&/      Meeting     ���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  �|W�,�  �(#&/      Meeting                        This_stuffs_This_stuffs_                                     Q�e�,�  r,#&/       Birthday U  p ��U  0��U  pSome_stuffs_Some_stuffs_ �U  0��U  ���U  p��U  0��U  ���,�  �S#&/      Some_stuffs                    Some_stuffs_Some_stuffs_                                     �c�#-�  0�-&/      Appointment ���U  ����U  0�Some_stuffs_Some_stuffs_ �U   ���U  ����U  ����U  @���U  ���#-�  ��-&/       Workout     P[��U  \��U  �`Some_stuffs_Some_stuffs_ �U   l��U  �l��U  �g��U  �h��U  ���#-�  z�-&/       Meeting     p���U  0���U  ��This_stuffs_This_stuffs_ �U  0���U  ����U  ����U  p���U  0�>$-�  ~$.&/       Meeting ffs ����U  p���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  �J$-�  �'.&/       Meeting     ����U  0���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �YK$-�  �'.&/      Workout     ����U  @���U   �Some_stuffs_Some_stuffs_ �U  @��U  ���U  @��U  ���U  B_L$-�  (.&/       Some_stuffs ���U  ���U  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  =��$-�  �H.&/      Birthday    ����U  @���U   �This_stuffs_This_stuffs_ �U   ���U  ����U  ����U  p���U  z�$-�  �M.&/       Workout ffs P-��U  �-��U  �.justforfun_justforfun_ _ �U  �0��U  �1��U   2��U  �2��U  `p�$-�  �O.&/       Birthday U  ����U   ���U  ��justforfun_justforfun_ ��U  @���U  ����U  @���U  ����U  �^%-�  Nn.&/      Appointment �9��U  �:��U  �>justforfun_justforfun_ ��U  0K��U  �K��U  �P��U  @Q��U  �l%-�  �q.&/       Some_stuffs ����U  `���U   �justforfun_justforfun_ ��U  `���U   ���U  ����U  ����U  �&�%-�  ��.&/       Birthday    ����U  P���U  �justforfun_justforfun_ ��U  ���U  ����U  ����U  ����U  �1&-�  k�.&/       Some_stuffs ����U  0���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  J&-�  ��.&/       Meeting     0���U   ���U  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `���U  |2&-�  ��.&/      Meeting �U   o��U  �o��U  �pjustforfun_justforfun_ ��U  Ps��U  t��U  �t��U  �u��U  ��&-�  �.&/      Birthday    ���U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ���&-�  y�.&/       Some_stuffs ����U  P���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �&-�  U�.&/       Workout     P=��U  >��U  �>This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  PC��U  9�.'-�  �.&/       Birthday                       Some_stuffs_Some_stuffs_                                     \e;'-�  K�.&/      Workout                        This_stuffs_This_stuffs_                                     �'-�  �/&/      Workout     P[��U  \��U  �`Some_stuffs_Some_stuffs_ �U   l��U  �l��U  �g��U  �h��U  ���'-�  �/&/       Workout     `f��U   g��U   lSome_stuffs_Some_stuffs_ �U  pj��U  0k��U  �q��U  �r��U  �9`(-�  B3/&/       Some_stuffs 0���U  ����U  p�This_stuffs_This_stuffs_ �U  P
��U  �
��U  @���U  ����U  �W{(-�  3:/&/      Birthday    �B��U  pC��U  0DThis_stuffs_This_stuffs_ �U  pF��U  0G��U  �G��U  0H��U  ��(-�  ?Z/&/       Birthday    `"��U  �"��U  `#Some_stuffs_Some_stuffs_ �U  �%��U   &��U  �&��U   '��U  ��)-�  �_/&/       Some_stuffs  ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `���U  R�)-�  �/&/       Appointment ����U  @���U  ЋSome_stuffs_Some_stuffs_ �U  ����U  `���U   ���U  ����U  �ޛ)-�  �/&/       Some_stuffs ���U  @��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  � ��U  $i�)-�  ��/&/      Meeting �U   ���U  ����U  ��justforfun_justforfun_ ��U  ����U  P���U  ���U  й��U  9�)-�  ��/&/       Some_stuffs 0f��U  �g��U  �iSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �t��U  ��1*-�  z�/&/       Meeting     ����U  ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `���U  �zB*-�  ��/&/       Some_stuffs �H��U  �I��U  0Jjustforfun_justforfun_ ��U  �L��U  �M��U  @^��U  �^��U  X��*-�  ��/&/       Appointment ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  ��*-�  ��/&/      Appointment 0f��U  �g��U  �iSome_stuffs_Some_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  �?\+-�  ��/&/       Birthday    ����U  `���U  ��This_stuffs_This_stuffs_ �U  ����U  `���U  е��U  ����U  c!c+-�  ��/&/       Birthday    �R��U  PS��U  TThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �W��U  Q�j+-�  ��/&/       Appointment ����U  P���U  �This_stuffs_This_stuffs_ �U  ����U  `���U  Э��U  P���U  ��w+-�  ��/&/      Birthday    ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  ���+-�  �0&/       Meeting     �]��U  @^��U  �^This_stuffs_This_stuffs_ �U  �`��U  �a��U  b��U  �b��U  <0,-�  �!0&/      Some_stuffs ���U  Ш��U  ��Some_stuffs_Some_stuffs_ �U  P���U  ���U  ����U  ���U  �V�,-�  �F0&/      Appointment ����U  `���U   �This_stuffs_This_stuffs_ �U  ����U  p���U  0���U  ����U   '<--�  �q0&/       Workout     0D��U  �D��U  0ESome_stuffs_Some_stuffs_ �U  �G��U  0H��U  �H��U  �I��U  X}�--�  G�0&/       Appointment 0f��U  �g��U  �ijustforfun_justforfun_ ��U  �p��U  �q��U  �s��U  �t��U  ��--�  ��0&/      Birthday    �]��U  �n��U  `_justforfun_justforfun_ ��U   b��U  �b��U   c��U  �c��U  2��--�  >�0&/       Some_stuffs                    justforfun_justforfun_                                       ̊b.-�  �0&/      Workout     ���U  ����U  P�Some_stuffs_Some_stuffs_ �U  @���U  ���U  ���U  ����U  ��.-�  ��0&/      Appointment @	��U  �	��U  @	This_stuffs_This_stuffs_ �U  �	��U  `		��U  �		��U  `
	��U  �M/-�  E�0&/       Meeting �U  0f��U  �g��U  �iThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �t��U  �N�/-�  �1&/      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_              ڗ/-�  @1&/       Birthday    ����U  0���U  ��justforfun_justforfun_ ��U  ����U  p���U  0���U  ���U  � �0-�  �V1&/      Appointment 0���U   ���U  @�This_stuffs_This_stuffs_ �U  p���U  0���U  ����U  `���U  ��0-�  vX1&/       Appointment ��	��U  `�	��U  �	This_stuffs_This_stuffs_ �U  �	��U  `�	��U  �	��U  `�	��U  ��P1-�  }1&/       Some_stuffs P���U  ����U  P�justforfun_justforfun_ ��U  ���U  ����U  P���U  ���U  <�a1-�  w�1&/      Meeting                        justforfun_justforfun_                                       �>i1-�  d�1&/       Some_stuffs p���U  0���U  ��This_stuffs_This_stuffs_ �U  p���U  ����U  ����U  0���U  �On1-�  ��1&/       Workout     `"��U  �"��U  `#This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   '��U  -�1-�  $�1&/      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �E�1-�  �1&/       Birthday nt `���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `���U  j�2-�  q�1&/       Appointment `���U  �.	��U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  }�2-�  ?�1&/      Appointment ����U  p���U  0�This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U   ���U  &�2-�  ��1&/       Workout �U  0���U   ���U  @�Some_stuffs_Some_stuffs_ �U  p���U  0���U  ����U  `���U  ��2-�  ��1&/       Meeting     @��U  ���U  @This_stuffs_This_stuffs_ �U  ���U  ���U   ��U  ���U  8d3-�  ��1&/      Some_stuffs 0f��U  �g��U  �ijustforfun_justforfun_ ��U  �p��U  �q��U  �s��U  �t��U  �,3-�  ��1&/       Workout �U  0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  �f3-�  ��1&/       Meeting �U  0f��U  �g��U  �iThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �t��U  PT$3-�  ��1&/       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ��)3-�  E�1&/       Workout                        This_stuffs_This_stuffs_                                     c303-�  ��1&/       Workout     е��U  ����U  �justforfun_justforfun_ ��U  ����U  ����U  ���U  ����U  �13-�  ?�1&/       Birthday    P���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �|63-�  x�1&/       Some_stuffs `���U   ���U  НSome_stuffs_Some_stuffs_ �U  0���U  ���U  ����U  p���U  �]�3-�  A2&/       Birthday                       justforfun_justforfun_                                       ���3-�  �2&/      Some_stuffs  ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  2u�3-�   2&/       Birthday    @���U  ����U  p�Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   ���U   �H4-�  �?2&/       Birthday    ����U  @���U  �Some_stuffs_Some_stuffs_ �U  P���U  ���U   ���U  ����U  �]L4-�  �@2&/      Appointment �9��U  �:��U  �>Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @Q��U  �ZS4-�  eB2&/       Appointment ����U  `���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  3�g4-�  �G2&/       Some_stuffs ���U  P��U  justforfun_justforfun_ ��U  P��U  ���U  P��U  ��U  p��4-�  &g2&/       Some_stuffs P���U  ���U  p�This_stuffs_This_stuffs_ �U  ����U  ����U  @���U    ��U  ��4-�  *g2&/       Birthday    p��U  ���U  �Some_stuffs_Some_stuffs_ �U  p"��U  �"��U  �#��U  p$��U  ��4-�  zi2&/      Birthday     ���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��4-�  �l2&/       Appointment `���U  ���U  ��Some_stuffs_Some_stuffs_ �U  ����U  ���U  ����U  ���U  �<_-�  �>=&/       Some_stuffs �8��U  p9��U  �9Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ?��U  �K_-�  �B=&/      Birthday U   ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  p���U  ���U  ж��U   w�_-�  �c=&/       Birthday    p;��U  �;��U  P=justforfun_justforfun_ ��U  �?��U  P@��U  A��U  �A��U  ���_-�  He=&/      Meeting     �6��U   7��U  �7Some_stuffs_Some_stuffs_ �U  P9��U  �9��U  p:��U  0;��U  j5�_-�  �e=&/       Birthday nt �k��U  `l��U   mSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �q��U  �=o`-�  �=&/      Appointment �b��U  @c��U  �cThis_stuffs_This_stuffs_ �U  �f��U  pg��U  0h��U  �h��U  ��a-�  e�=&/       Meeting     �d��U  �e��U  @fSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @j��U  �a-�  ��=&/      Appointment �	��U  0
��U  �
Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  ���U  }��a-�  ?�=&/      Some_stuffs  b��U  �b��U   cSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �g��U  �G�a-�  ��=&/       Some_stuffs  2��U  �2��U   3Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   7��U  ��a-�  ��=&/       Meeting     ���U  ����U  P�This_stuffs_This_stuffs_ �U  @���U  ���U  ���U  ����U  �'9b-�  X>&/       Workout      ���U  ����U  `�Some_stuffs_Some_stuffs_ �U   ���U  ����U  `���U   ���U  �:b-�  �>&/       Meeting     ����U  P���U  �justforfun_justforfun_ ��U  P���U  ����U  ����U  P���U  f�@b-�  @>&/      Birthday     ���U  ����U  0�This_stuffs_This_stuffs_ �U  0���U  ����U  ����U  p���U  p��b-�  �+>&/       Birthday nt ����U  0���U  �This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  0���U  8R|c-�  U>&/       Workout     �C��U  �D��U  @ESome_stuffs_Some_stuffs_ �U  �G��U   H��U  �H��U  @I��U  "yd-�  �x>&/       Workout     �}��U  p~��U  �~This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Ђ��U  y�d-�  �y>&/       Workout ffs ����U  p���U  0�justforfun_justforfun_ ��U  ����U  0���U  P
��U  �
��U  p d-�  �{>&/       Workout     `V��U   W��U  �WThis_stuffs_This_stuffs_ �U  �Z��U  �[��U  @\��U   ]��U  �Ѡd-�  ��>&/      Meeting �U  0f��U  �g��U  �iSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �t��U  "Ţd-�  t�>&/       Workout     м��U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  	�d-�  �>&/       Birthday U  ����U  p���U  ��justforfun_justforfun_ ��U  ����U  p���U  ����U  p���U  1-*e-�  �>&/       Workout  fs P���U  ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  @�0e-�  ��>&/       Appointment �o��U   p��U  �pjustforfun_justforfun_ ��U   s��U  �s��U   t��U  �t��U  ��e-�  ��>&/       Workout     ����U  @���U   �This_stuffs_This_stuffs_ �U  ���U  ж��U  ����U  P���U  ��^f-�  -?&/       Some_stuffs P���U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  1<`f-�  ~?&/       Some_stuffs 0f��U  �g��U  �iSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �t��U  3�af-�  �?&/       Some_stuffs ���U  ����U  ��justforfun_justforfun_ ��U  ����U  @���U  0���U   ���U  H�df-�  �?&/       Appointment ����U  `���U  ��This_stuffs_This_stuffs_ �U  ����U  `���U  е��U  ����U  �!�f-�  �7?&/       Meeting     p��U  ���U  �Some_stuffs_Some_stuffs_ �U  p"��U  �"��U  �#��U  p$��U  `-�f-�  8?&/       Birthday     ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  `���U   ���U  ����U  ��g-�  ??&/      Meeting     ��U  ���U  PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �	��U  BI�g-�  H^?&/       Meeting     �}��U  `~��U   Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `���U  ��g-�  �a?&/      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �5�g-�  ne?&/       Meeting      W��U  �W��U  @Xjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  �\��U  ~�3h-�  �?&/      Workout      V��U  �V��U  �WThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0[��U  ��3h-�  +�?&/       Workout     0���U  ����U  ��Some_stuffs_Some_stuffs_ �U  p���U  0���U  ����U  ����U  ��3h-�  +�?&/       Appointment ���U  0 ��U  � Some_stuffs_Some_stuffs_ �U  �#��U  p$��U  0%��U  �3��U  %��h-�  ��?&/      Some_stuffs @��U  ���U  @This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  l�h-�  U�?&/       Workout     0���U  ���U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��_i-�  ��?&/      Appointment 0���U   ���U  @�Some_stuffs_Some_stuffs_ �U  p���U  0���U  ����U  `���U  Rqgi-�  ��?&/       Some_stuffs @�	��U  �	��U  p�	Some_stuffs_Some_stuffs_ �U  ��	��U  `�	��U  ��	��U  `�	��U  3�mi-�  ��?&/       Birthday    `��U   ��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �!��U  �1oi-�  ��?&/       Some_stuffs 0���U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  q��i-�  ��?&/       Workout     ��U  ���U  �Some_stuffs_Some_stuffs_ �U  ���U  ���U  p��U  0��U  J�j-�  }@&/       Some_stuffs ���U  0��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0��U  ,hj-�  -@&/      Meeting     ����U  @���U  P�This_stuffs_This_stuffs_ �U  P���U  Т��U  ����U  P���U  �ٟj-�  �(@&/       Some_stuffs @��U  ���U  @Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �ˤj-�  0*@&/       Workout     0���U  ���U  ��This_stuffs_This_stuffs_ �U  ����U  0���U  ���U  p���U  D9"k-�  LJ@&/      Birthday    ����U  @���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �,�k-�  �o@&/      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �_�k-�  r@&/       Meeting  U   ���U  ����U   �justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ���U  q�k-�  Fv@&/       Appointment ���U  ����U  0�Some_stuffs_Some_stuffs_ �U   ���U  ����U  ����U  @���U  �pl-�  @&/       Appointment ���U  ж��U  ��Some_stuffs_Some_stuffs_ �U  P���U  ���U  л��U  ����U  @C�l-�  ��@&/       Birthday    �`��U  �a��U  `fjustforfun_justforfun_ ��U  �g��U  �h��U  pj��U  0k��U  �l-�  9�@&/      Birthday    �^��U  @_��U  �_This_stuffs_This_stuffs_ �U  @b��U  �b��U  �c��U  @d��U  ��m-�  ��@&/      Some_stuffs  b��U  �b��U   cThis_stuffs_This_stuffs_ �U  �e��U  `f��U  �f��U  �g��U  A��m-�  �@&/       Appointment ����U   ���U  ��justforfun_justforfun_ ��U  ���U  ����U  ���U  ����U  y%n-�  �A&/       Meeting �U  0f��U  �g��U  �ijustforfun_justforfun_ ��U  �p��U  �q��U  �s��U  �t��U  01n-�  �A&/       Workout     p��U  0��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  x�n-�  �5A&/       Appointment                    This_stuffs_This_stuffs_                                     �@�n-�  �5A&/      Birthday fs p���U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  b�Io-�  �ZA&/       Appointment @'��U   (��U  �(This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �-��U  �
Ko-�  �ZA&/       Meeting     ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��Ro-�  �\A&/       Workout �U  0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  ��do-�  �aA&/      Workout     P���U  ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  �;�o-�  ځA&/       Birthday U  ����U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  p���U  0���U  ����U  ���o-�  ��A&/       Appointment  h��U  �h��U   ijustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  �m��U  ���o-�  Z�A&/       Appointment `���U   ���U  ��Some_stuffs_Some_stuffs_ �U  ����U  `���U   ���U  ����U  :l p-�  S�A&/       Meeting     0U��U  �U��U  `VThis_stuffs_This_stuffs_ �U  @Y��U   Z��U  �Z��U  �[��U  `*yp-�  <�A&/       Birthday                       justforfun_justforfun_                                       ��p-�  ��A&/      Meeting      ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  )�p-�  �A&/       Some_stuffs p��U  0��U  0This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p0��U  ���p-�  C�A&/       Some_stuffs 0"��U  �<��U  0$justforfun_justforfun_ ��U  �&��U  �'��U  0(��U  �(��U  �q-�  ��A&/      Birthday    ��U  ���U  �This_stuffs_This_stuffs_ �U  ���U  ���U  p��U  0��U  �'q-�  ��A&/       Some_stuffs 0���U  ����U  p�justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  ����U  YQ˚-�  �}L&/       Workout     е��U  ����U  �Some_stuffs_Some_stuffs_ �U  ����U  ����U  ���U  ����U  �W՚-�  X�L&/       Workout     �+��U  �,��U  P-justforfun_justforfun_ ��U  �/��U  `0��U  �0��U  �1��U  �'�-�  /�L&/      Meeting     ����U  p���U  0�Some_stuffs_Some_stuffs_ �U  ����U  ����U  p ��U  0��U  ��{�-�  ��L&/       Appointment �h	��U  `i	��U  j	This_stuffs_This_stuffs_ �U  l	��U  �l	��U  @m	��U  �m	��U  D��-�  ��L&/      Appointment �t��U  �u��U  vSome_stuffs_Some_stuffs_ �U  `y��U   z��U  �z��U  `{��U  ���-�  ��L&/       Workout  U  0f��U  �g��U  �iSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  �t��U  X�	�-�  G�L&/       Birthday                       This_stuffs_This_stuffs_                                     �$�-�  ��L&/      Birthday    p�	��U   �	��U  ��	justforfun_justforfun_ 	��U  ��	��U  `�	��U  ��	��U  `�	��U  X/��-�  ��L&/       Meeting �U   ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �.��-�  �L&/      Workout     @���U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  �/�-�  eM&/       Meeting     p ��U  0��U  pSome_stuffs_Some_stuffs_ �U  0��U  ���U  p��U  0��U  �VA�-�  M&/      Meeting ffs �/��U  p0��U  �4Some_stuffs_Some_stuffs_ �U  �>��U  �?��U   E��U  �F��U  �J�-�  N!M&/       Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             c+P�-�  �"M&/       Appointment 0��U  ���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0 ��U  ��˝-�  �BM&/       Workout �U  � ��U  �!��U  p"This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   (��U  "�-�  @IM&/       Some_stuffs ����U  @���U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  z�-�  {IM&/       Meeting     ����U  P���U  ��This_stuffs_This_stuffs_ �U   ���U  ����U   ���U  ����U  ��g�-�  ejM&/       Meeting �U  ����U  0���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  1�m�-�  �kM&/       Appointment p:��U  0;��U  �;Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �?��U  o�-�  NlM&/      Appointment  ]	��U  �]	��U   ^	Some_stuffs_Some_stuffs_ �U   `	��U  �`	��U   a	��U  �a	��U  �;~�-�  0pM&/       Some_stuffs  ���U  ����U  `�This_stuffs_This_stuffs_ �U  ����U  ���U  ����U  ���U  ��-�  d�M&/      Appointment л��U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  aK�-�  ܖM&/       Workout     `���U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  P��-�  �M&/       Meeting      o��U  �o��U  �pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �u��U  \�)�-�  ��M&/      Meeting �U  p��U  0��U  0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p0��U  �q/�-�  �M&/       Birthday nt 0���U  ����U  p�This_stuffs_This_stuffs_ �U  ����U  0���U  ���U  p���U  ��@�-�  ��M&/       Some_stuffs 05��U  �5��U  06This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �:��U  �XǠ-�  �N&/       Appointment `���U   ���U  НThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  D�Π-�  �N&/      Birthday                       Some_stuffs_Some_stuffs_                                     rp�-�  D1N&/      Birthday    @���U  ����U  ��This_stuffs_This_stuffs_ �U   ���U  ����U  @���U  ����U  )�-�  IVN&/       Some_stuffs  a��U  �a��U  @bThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �f��U  ,"�-�  m[N&/      Appointment � ��U  �!��U  p"Some_stuffs_Some_stuffs_ �U  0%��U  �3��U  @'��U   (��U  �鐢-�  {N&/      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             @MC�-�  ȨN&/       Some_stuffs ����U  ����U  �This_stuffs_This_stuffs_ �U  ����U  `���U  @���U  ���U   "£-�  @�N&/       Workout ent �/��U  p0��U  �4Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �F��U  <e�-�  ��N&/      Some_stuffs  ��U  ���U   This_stuffs_This_stuffs_ �U  `��U  ���U  `��U   ��U  �_�-�  �O&/      Meeting      ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ���-�  �=O&/       Birthday nt  ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  `���U  ����U  `���U  ����-�  c@O&/       Appointment �t��U  �u��U  vSome_stuffs_Some_stuffs_ �U  `y��U   z��U  �z��U  `{��U  = ��-�  �CO&/      Appointment p���U  ����U  p�This_stuffs_This_stuffs_ �U  ����U  ����U   ���U  ����U  �#�-�  _eO&/       Appointment 00��U  �0��U  p1Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �5��U  t=5�-�  �iO&/      Workout     0���U  ����U  p�Some_stuffs_Some_stuffs_ �U  ����U   ���U  @���U   ���U   �˦-�  `�O&/       Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             S7ͦ-�  ��O&/       Some_stuffs 0���U  ����U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  )Oئ-�  ��O&/       Birthday U   b��U  �b��U   cThis_stuffs_This_stuffs_ �U  �e��U  `f��U  �f��U  �g��U  ��٦-�  �O&/      Appointment �}��U  p~��U  �~Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  Ђ��U  I�V�-�  ݳO&/       Workout     pv��U  0w��U  �wSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0|��U  R0`�-�  R�O&/       Some_stuffs  ���U  ����U  `�Some_stuffs_Some_stuffs_ �U   ���U  ����U  `���U   ���U  ��p�-�  ��O&/      Some_stuffs �<��U  �=��U   >This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �A��U  �-�  ��O&/      Workout     �Z��U  �[��U  @\This_stuffs_This_stuffs_ �U  `_��U   `��U  �`��U  `a��U  �0�-�  ��O&/       Appointment �K��U  0L��U  �LThis_stuffs_This_stuffs_ �U  �O��U  pP��U  �P��U  �Q��U  <q��-�  wP&/      Workout ffs @X��U  �X��U  �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ^��U  ��*�-�  �+P&/       Some_stuffs ����U  p���U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  a�/�-�  �,P&/       Appointment  ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  0��U  ����U  p���U  jK:�-�  �/P&/       Appointment P9��U  �9��U  p:Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �>��U  ©-�  uRP&/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��ө-�  �VP&/       Some_stuffs @T��U  �T��U  @Ujustforfun_justforfun_ ��U  �W��U  @X��U  �X��U  @Y��U  �qK�-�  �uP&/      Workout     P���U  Є��U  ��This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  ����U  �n[�-�  �yP&/       Some_stuffs ����U  `���U   �This_stuffs_This_stuffs_ �U  ����U  `���U  ����U  `���U  ^�-�  _zP&/       Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             L�-�  �P&/      Appointment �P��U  �Q��U  pRjustforfun_justforfun_ ��U  0U��U  �U��U  `V��U   W��U  A+�-�  ��P&/       Workout     ����U  ����U  P�This_stuffs_This_stuffs_ �U  ���U  ����U  ����U  P���U  "$��-�  ԡP&/       Some_stuffs `���U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  mD��-�  U�P&/      Appointment p���U  ���U  ��Some_stuffs_Some_stuffs_ �U  ���U  ж��U  P���U  ���U  b֛�-�  ��P&/       Workout ent  +��U  �+��U  �/This_stuffs_This_stuffs_ �U  �9��U  �:��U  �>��U  �?��U  ���-�  �P&/       Workout     ����U  `���U  ��justforfun_justforfun_ ��U  ����U  `���U  е��U  ����U  ���-�  k�P&/       Workout ffs ����U  ����U  `�justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ���U  ���-�  ~�P&/      Meeting �U  �
��U  ���U  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0��U  �k�-�  j�[&/       Appointment 0��U  ���U  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �"��U  �$x�-�  ��[&/       Workout     p��U  ���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �|�-�  ��[&/      Some_stuffs ���U  p��U  0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ���-�  x�[&/       Some_stuffs  ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  `���U  ����U  `���U  в��-�  ��[&/       Meeting     ���U  P��U   Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �y�-�  ��[&/      Meeting     P���U  ���U  лjustforfun_justforfun_ ��U  ���U  ����U  0���U  ���U  侞�-�  \&/      Meeting �U   ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �/�-�  95\&/      Meeting �U  P���U  ����U  P�This_stuffs_This_stuffs_ �U  ����U  P���U  ���U  ����U  (|��-�  �a\&/       Some_stuffs P���U  ����U  P�This_stuffs_This_stuffs_ �U  ����U  P���U  ����U  ����U  ��i�-�  ��\&/       Birthday    е��U  ����U  �This_stuffs_This_stuffs_ �U  ����U  ����U  ���U  ����U  $Em�-�  x�\&/      Some_stuffs ����U  p���U  0�Some_stuffs_Some_stuffs_ �U  ����U  0���U  ���U  ����U  ����-�  �\&/       Birthday     ���U  ����U  ��justforfun_justforfun_ ��U  Н��U  ����U  ����U  p���U  ��-�   �\&/       Meeting     ����U  p���U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  Bc�-�  ��\&/       Meeting ffs ����U  p���U  Љjustforfun_justforfun_ _ �U  ���U  ����U  ���U  ����U  �*�-�  >�\&/      Workout �U  ����U  @���U  �justforfun_justforfun_ ��U  P���U  ���U   ���U  ����U  h���-�  �\&/       Workout ent �'��U  P(��U  �(This_stuffs_This_stuffs_ �U  �*��U  P+��U  �+��U  �,��U  �׫�-�  �\&/      Meeting     �+��U   ,��U  �,Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �1��U  j9�-�  D�\&/      Birthday    p-��U  0.��U  �.This_stuffs_This_stuffs_ �U  p1��U  �1��U  �2��U  p3��U  *A�-�  @�\&/       Workout     �P��U  Q��U  �QSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �U��U  ��K�-�  � ]&/       Some_stuffs ����U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ���-�  , ]&/       Birthday    ���U  `��U  Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ���U  L3��-�  a#]&/      Birthday    ����U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ipd�-�  �H]&/       Appointment ����U  0���U  ��Some_stuffs_Some_stuffs_ �U  ����U  p���U  0���U  ���U  x�s�-�  �L]&/       Birthday    0r��U  �r��U  �sThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  px��U  ����-�  n]&/      Birthday    ����U  ����U   �Some_stuffs_Some_stuffs_ �U   ���U  ����U   ���U  ����U  �q �-�  �p]&/       Birthday fs  -��U  �-��U   .This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U   2��U  ꥞�-�  A�]&/       Some_stuffs @���U   ���U  ��justforfun_justforfun_ _ �U  ����U  @���U   ���U  p���U  ���-�  ��]&/      Birthday    �C��U  �D��U  EThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  I��U  1.��-�  ��]&/       Workout ffs  ���U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  K%�-�  ��]&/      Meeting     е��U  ����U  �This_stuffs_This_stuffs_ �U  ����U  ����U  ���U  ����U  ɻ4�-�  ��]&/       Some_stuffs �s	��U   t	��U  �t	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `x	��U  $��-�  �]&/      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             )(��-�  )�]&/       Appointment �8��U  p9��U  �9Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ?��U  �V�-�  �	^&/       Birthday    �]��U  @^��U  �^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �b��U  1i�-�  �^&/       Birthday                       justforfun_justforfun_ _                                     ��v�-�  ^&/      Workout �U  0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  ���-�  s2^&/      Some_stuffs  ��U  ���U  `oSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pt��U  P���-�  �W^&/       Birthday    �+��U   ,��U  �,This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �1��U  �%�-�  B�^&/       Birthday U  @���U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  <T%�-�  W�^&/      Some_stuffs ����U  ����U  p�Some_stuffs_Some_stuffs_ �U  0���U  ����U  ���U  ����U  Q�=�-�  ��^&/       Appointment  V��U  �V��U  �WThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  0[��U  Ec��-�  ��^&/      Meeting �U  0���U   ���U  @�Some_stuffs_Some_stuffs_ �U  p���U  0���U  ����U  `���U   ��-�  �^&/       Some_stuffs 0f��U  �g��U  �iThis_stuffs_This_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  �S�-�  ��^&/       Some_stuffs PL��U  M��U  �Mjustforfun_justforfun_ ��U  �P��U  Q��U  �Q��U  PR��U  �HS�-�  ��^&/       Birthday nt �{��U  0|��U  �|justforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U   ���U  �Bn�-�  ��^&/       Appointment Т��U  P���U  �Some_stuffs_Some_stuffs_ �U  Ц��U  ����U  ���U  Ш��U  ��r�-�  ��^&/       Meeting �U  е��U  ����U  �This_stuffs_This_stuffs_ �U  ����U  ����U  ���U  ����U  ,#t�-�  �^&/      Birthday                       Some_stuffs_Some_stuffs_                                     ���-�  �^&/       Workout      ��U  ���U  �This_stuffs_This_stuffs_ �U  0��U  ���U   $��U  �%��U  (��-�  ��^&/       Some_stuffs �t��U  �u��U  vSome_stuffs_Some_stuffs_ �U  `y��U   z��U  �z��U  `{��U  $���-�  �_&/      Workout                        Some_stuffs_Some_stuffs_                                     z��-�  �_&/       Birthday     4��U  �4��U  `5Some_stuffs_Some_stuffs_ �U  �7��U  `8��U   9��U  �9��U  �J��-�  a"_&/       Birthday    ����U  `���U  ��Some_stuffs_Some_stuffs_ �U  ����U  `���U  е��U  ����U  U)�-�  �E_&/      Appointment ���U  ����U  0�justforfun_justforfun_ ��U   ���U  ����U  ����U  @���U  ���-�  Xi_&/       Birthday     ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ዾ�-�  ,l_&/       Workout     �t��U  �u��U  vThis_stuffs_This_stuffs_ �U  `y��U   z��U  �z��U  `{��U  N��-�  !p_&/      Birthday    @���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  �Mf�-�  �_&/      Meeting     0���U  ����U  p�This_stuffs_This_stuffs_ �U  ����U   ���U  @���U   ���U  �u��-�  p�_&/       Meeting ent po	��U  �o	��U  pp	This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U   t	��U  l���-�  չ_&/      Workout     � ��U  �!��U  p"justforfun_justforfun_ ��U  0%��U  �3��U  @'��U   (��U  z�-�  �_&/      Some_stuffs                    justforfun_justforfun_                                       A��-�  ��_&/       Workout     p"��U  �"��U  �#Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �)��U  C�"�-�  �`&/       Some_stuffs ����U  `���U  ��justforfun_justforfun_ ��U   ���U  ����U   ���U  ����U  A�+�-�  (`&/       Birthday    0���U  ����U  0�This_stuffs_This_stuffs_ �U  p���U  0���U  ����U  0���U  �/�-�  	`&/      Birthday    ����U  @���U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  ��2�-�  `&/       Birthday    ���U  P���U  �Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  ���U  �}��-�  A0`&/       Workout     Р��U  ����U  P�This_stuffs_This_stuffs_ �U  ���U  ����U  ���U  ����U  ����-�  g1`&/      Birthday                       justforfun_justforfun_                                       �I�-�  =T`&/      Appointment ����U  ���U  ЮSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  0SS�-�  �V`&/       Workout                        justforfun_justforfun_                                       ��.�  Zk&/      Meeting     ����U  0���U  ��Some_stuffs_Some_stuffs_ �U  ����U  0���U  ����U  ����U  ��.�  �,k&/      Meeting ffs ���U  p���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  (�.�  �1k&/       Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             dj1.�  <Pk&/       Birthday nt @���U  ����U  `�justforfun_justforfun_ _ �U  `���U  ����U  ����U   ���U  V�4.�  Qk&/      Birthday U  �B��U  PC��U  �CThis_stuffs_This_stuffs_ �U  PF��U  �F��U  PG��U  �G��U  �k6.�  �Qk&/       Meeting     0���U   ���U  @�Some_stuffs_Some_stuffs_ �U  p���U  0���U  ����U  `���U  s�I.�  �Vk&/       Some_stuffs ����U  � ��U  @Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  �mQ.�  nXk&/       Workout     ����U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��.�  �wk&/       Appointment ����U   ���U  @�justforfun_justforfun_ ��U  @���U   ���U  ����U  @���U  �K�.�  �yk&/       Some_stuffs 0f��U  �g��U  �iThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �t��U  P�v.�  ��k&/       Some_stuffs �2��U  p3��U  04justforfun_justforfun_ ��U  06��U  �6��U  p7��U  08��U  �y.�  D�k&/      Meeting     ���U  ` ��U   !This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   %��U  �C.�  ��k&/       Birthday    �l��U  `m��U   justforfun_justforfun_ ��U  �p��U  �q��U  0r��U  �r��U  M=.�  ��k&/      Some_stuffs PO��U  �O��U  �PSome_stuffs_Some_stuffs_ �U  �R��U  PS��U  T��U  �T��U  ��.�  ��k&/       Workout     �Q	��U  R	��U  �R	justforfun_justforfun_ 	��U  �T	��U  @U	��U  �U	��U  @V	��U  !c�.�  4�k&/       Meeting     ���U   ��U  �Some_stuffs_Some_stuffs_ �U  p��U  ���U  ���U  @��U  p�.�  ��k&/      Appointment ����U  @���U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  P�C.�  �l&/       Birthday    ����U  @���U  �This_stuffs_This_stuffs_ �U  P���U  ���U   ���U  ����U  �jF.�  8l&/       Birthday     ���U  ����U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  ��L.�  �l&/      Birthday nt ����U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  ��.�  �:l&/       Meeting     0"��U  �<��U  0$justforfun_justforfun_ ��U  �&��U  �'��U  0(��U  �(��U  ��.�  �=l&/       Workout     �B��U  pC��U  �CSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   H��U  �/�.�  �Bl&/      Appointment ����U  0���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �0g.�  %dl&/       Appointment  !��U  �!��U  `"Some_stuffs_Some_stuffs_ �U  �$��U   %��U  �%��U   &��U  \�k.�  Kel&/      Workout �U  0f��U  �g��U  �iSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �t��U  �Wt.�  �gl&/       Meeting     �<��U  �=��U   >justforfun_justforfun_ _ �U  �N��U  PO��U  0A��U  �A��U  ��.�  �jl&/       Some_stuffs ����U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  ��.�  �jl&/       Meeting     `���U  ����U  `�justforfun_justforfun_ ��U  ����U  `���U   ���U  ����U  ��.�  Z�l&/      Some_stuffs @(��U  �(��U  p)This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  �-��U  ��.�  o�l&/       Workout                        This_stuffs_This_stuffs_                                     �Ǯ.�  �l&/       Birthday    ���U  @	��U  �	justforfun_justforfun_ _ �U   ��U  ���U  @��U  ���U  ,X0.�  -�l&/      Some_stuffs ����U  0���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  �=5.�  n�l&/       Birthday fs Pb	��U  �b	��U  Pc	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `g	��U  ��B.�  ��l&/       Appointment ����U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  Q��.�  ��l&/       Workout      ���U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  t��.�  jm&/      Appointment �z��U  `{��U   |This_stuffs_This_stuffs_ �U  p��U  0���U  ����U  ����U  T�f.�  �(m&/      Meeting     ����U  p���U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �r.�  �+m&/       Workout     ����U  @���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �_�.�  -Nm&/       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ���.�  �Om&/      Meeting     �t��U  �u��U  vSome_stuffs_Some_stuffs_ �U  `y��U   z��U  �z��U  `{��U  �q.�  �Pm&/       Some_stuffs                    Some_stuffs_Some_stuffs_                                     �^�.�  tm&/       Some_stuffs �f��U  �g��U  `hThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `m��U  ��".�  P�m&/       Meeting     Н��U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  @ $.�  ��m&/       Appointment  o��U  �o��U  �pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �u��U  1L+.�  ~�m&/       Meeting     0r��U  �r��U  �sThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  px��U  �?.�  ��m&/      Workout �U  ��	��U  @�	��U  ��	justforfun_justforfun_ 	��U  ��	��U  p�	��U  ��	��U  p�	��U  )��.�  I�m&/       Workout     p ��U  0��U  pSome_stuffs_Some_stuffs_ �U  0��U  ���U  p��U  0��U  $��.�  X�m&/      Some_stuffs                    Some_stuffs_Some_stuffs_                                     Q,a.�  ��m&/       Workout      ���U  ����U  ��justforfun_justforfun_ ��U  ����U  `���U   ���U  ����U  ފl.�  ��m&/      Birthday    ����U  ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  Ёr.�  B�m&/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �r�.�  �n&/      Appointment �p��U  �q��U  0rThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0w��U  8��.�  Sn&/       Birthday    ����U  0���U  ��Some_stuffs_Some_stuffs_ �U  @���U  ����U  @���U  ����U  ��.�  �6n&/      Birthday nt 0f��U  �g��U  �iSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �t��U  �a�.�  k8n&/       Appointment 0���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��.�  p<n&/       Workout     �B��U  pC��U  0DSome_stuffs_Some_stuffs_ �U  pF��U  0G��U  �G��U  0H��U  � .�  :^n&/      Meeting                        This_stuffs_This_stuffs_                                     1�4.�  ~cn&/       Meeting      ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ж��U  X�.�  �n&/       Birthday    ����U  `���U  ��Some_stuffs_Some_stuffs_ �U  ����U  `���U  е��U  ����U  ��.�  s�n&/      Some_stuffs �C��U  �D��U  @Ejustforfun_justforfun_ _ �U  �G��U   H��U  �H��U  @I��U  Z��.�  ��n&/       Workout ffs ����U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0��U  ��.�  �n&/       Workout     ����U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ô�.�  x�n&/       Some_stuffs  ���U  ����U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  hzk .�  �n&/       Meeting �U  0���U  ����U  p�justforfun_justforfun_ ��U  ����U   ���U  @���U   ���U  7�� .�  ~�n&/       Birthday fs �l��U  `m��U   This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �r��U  TB� .�  ��n&/       Birthday    Ъ��U  ����U  P�justforfun_justforfun_ _ �U  Ю��U  ����U  ���U  ����U  :.� .�  ��n&/       Appointment  ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  �Z� .�  ��n&/      Appointment ����U  `���U   �This_stuffs_This_stuffs_ �U   ���U  ����U  ����U  `���U  c�!.�  |�n&/       Workout     ���U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��!.�  ��n&/       Meeting     ����U  ����U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  UA!.�  ��n&/       Meeting     �H��U  @I��U  �Ijustforfun_justforfun_ ��U  �K��U  @L��U  �L��U  �M��U  ��!.�  Z�n&/       Appointment �'��U  P(��U  �(Some_stuffs_Some_stuffs_ �U  �*��U  P+��U  �+��U  �,��U  �N�!.�  ��n&/       Workout     ����U  @���U   �Some_stuffs_Some_stuffs_ �U  ���U  ж��U  ����U  P���U  �!.�  5�n&/       Appointment �X��U  Y��U  �YThis_stuffs_This_stuffs_ �U  �[��U  `\��U  �\��U  `]��U  �:�!.�   o&/       Birthday    ���U  ����U  0�This_stuffs_This_stuffs_ �U   ���U  ����U  ����U  @���U  ���!.�  so&/      Some_stuffs `���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `���U  �Y$".�  �#o&/       Meeting ffs  ���U  ����U  ��Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  p���U  ��0".�  'o&/       Birthday    `o��U   p��U  �pThis_stuffs_This_stuffs_ �U  �s��U  pt��U  0u��U  �u��U  I"�".�  �Ho&/       Appointment  5��U  �5��U  �6This_stuffs_This_stuffs_ �U  �_��U  @`��U  P9��U  �9��U  N��".�  aIo&/      Workout ffs ���U  ����U  p�justforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U  P���U  ���".�  �Ko&/       Workout ffs  5��U  �5��U  �6justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  �9��U  mI#.�  �no&/       Appointment `���U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  %Z#.�  8so&/      Birthday    Т��U  P���U  �Some_stuffs_Some_stuffs_ �U  Ц��U  ����U  ���U  Ш��U  5b�#.�  B�o&/      Meeting     0���U  ����U  ��justforfun_justforfun_ ��U  p���U  0���U  ����U  ����U   ��#.�  ��o&/       Meeting     ����U  ���U  гSome_stuffs_Some_stuffs_ �U  ����U  0���U  ����U  p���U  I�M.�  �Ez&/       Some_stuffs ����U  0���U  ��This_stuffs_This_stuffs_ �U  ����U  p���U  0���U  ����U  l¡M.�  Fz&/      Appointment ��U  ���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0��U  b/�M.�  \Mz&/       Appointment  g��U  �g��U   hSome_stuffs_Some_stuffs_ �U  �j��U  `k��U  �k��U  `l��U  ���N.�  :�z&/       Some_stuffs 0>��U  �>��U  p?This_stuffs_This_stuffs_ �U  pA��U  �A��U  pB��U  �B��U  ��N.�  ��z&/      Some_stuffs P���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  |�uO.�  ߽z&/      Appointment p��U  0��U  �Some_stuffs_Some_stuffs_ �U  �	��U  0
��U  �
��U  ���U  R�uO.�  �z&/       Meeting     ���U  ����U  ��justforfun_justforfun_ ��U  ����U  @���U  0���U   ���U  �G�O.�  Z�z&/       Workout     �L��U  �M��U  @^This_stuffs_This_stuffs_ �U  �P��U  �Q��U  pR��U  �R��U  t��P.�  j
{&/      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             r��P.�  �{&/       Meeting ent @��U  ���U  ��This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  )��P.�  	{&/       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �)9Q.�  s1{&/      Birthday    �K��U  0L��U  �LThis_stuffs_This_stuffs_ �U  �O��U  pP��U  �P��U  �Q��U  !&OQ.�  7{&/       Birthday    @E��U  �E��U  �Fjustforfun_justforfun_ ��U  �H��U  @I��U  �I��U  @J��U  �8�Q.�  y\{&/       Meeting     p���U  ����U  ��Some_stuffs_Some_stuffs_ �U  @���U  ����U  ����U   ���U  ���Q.�  /^{&/      Workout                        This_stuffs_This_stuffs_                                     aR.�  5}{&/       Meeting                        This_stuffs_This_stuffs_                                     �FlR.�  �{&/      Meeting ffs `���U  ����U  ��justforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U  P���U  �NuR.�  b�{&/       Some_stuffs ��U  ���U  PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �	��U  ��R.�  �{&/       Workout     ���U  p��U  0This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  ���U  �l�R.�  |�{&/      Workout ffs ���U  Ѓ��U  ��justforfun_justforfun_ _ �U  ���U  ����U  P���U  Ј��U  F S.�  ��{&/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �S.�  է{&/       Workout     ���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  I�S.�  ��{&/       Meeting     0��U  ���U  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0
��U  �`S.�  !�{&/       Workout     �,��U  �-��U  @.This_stuffs_This_stuffs_ �U   1��U  �1��U  �2��U   3��U  �S.�  6�{&/       Meeting      o��U  �o��U  �pSome_stuffs_Some_stuffs_ �U  Ps��U  t��U  �t��U  �u��U  ly�S.�  u�{&/      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �6T.�  G�{&/      Workout     ����U  p���U  0�Some_stuffs_Some_stuffs_ �U  ���U  ����U  p���U  ����U  ���T.�  �|&/       Meeting     ���U  @��U  �justforfun_justforfun_ ��U  0��U  ���U  0E��U  �E��U  �%�T.�  n|&/       Birthday    �L��U  �M��U  @NThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   R��U  ���T.�  �|&/       Birthday nt ����U  `���U  ��Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ����U  ���T.�  ~ |&/      Meeting                        justforfun_justforfun_                                       tI�U.�  Ji|&/      Birthday     ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ж��U  �B�U.�  j|&/       Birthday    0��U  ���U  �This_stuffs_This_stuffs_ �U  0��U  ���U  ���U  0 ��U  P��V.�  ��|&/       Birthday    ���U  ����U  P�This_stuffs_This_stuffs_ �U  ���U  Ш��U  ����U  P���U  Ai�V.�  H�|&/       Appointment ����U  `���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �ťV.�  �|&/      Meeting     ����U  @���U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  ���V.�  d�|&/       Meeting     �S��U  pT��U  0USome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   Z��U  T�3W.�  V�|&/      Appointment                    justforfun_justforfun_                                       D�W.�  l�|&/      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             y"�W.�  ��|&/       Birthday     ���U  ����U  @�This_stuffs_This_stuffs_ �U  @���U  ����U  ����U   ���U  �hhX.�  L}&/       Meeting     0���U  ���U  ��Some_stuffs_Some_stuffs_ �U  ����U  0���U  ���U  p���U  � mX.�  y	}&/       Birthday    �W��U  �X��U  @Yjustforfun_justforfun_ ��U  @\��U   ]��U  �]��U  �n��U  �&wX.�  }&/      Some_stuffs pr��U  �r��U  �sSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �w��U  |k�X.�  _+}&/      Birthday    е��U  ����U  �Some_stuffs_Some_stuffs_ �U  ����U  ����U  ���U  ����U  �� Y.�  E/}&/       Some_stuffs  u��U  �u��U   vSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  z��U  وY.�  #R}&/      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��1Z.�  m}}&/       Meeting     0K��U  �K��U  �PSome_stuffs_Some_stuffs_ �U  P[��U  \��U  �`��U  �a��U  U�BZ.�  ��}&/      Meeting     0���U  ����U  �justforfun_justforfun_ ��U  p���U  ����U  p���U  0���U  ���Z.�  N�}&/       Birthday    ����U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  AY�Z.�  H�}&/       Meeting     �u��U  v��U  �vThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P{��U  ٓV[.�  W�}&/       Birthday    0���U   ���U  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `���U  *QX[.�  ��}&/       Appointment `k��U   l��U  �lSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �q��U  4�`[.�  ��}&/      Workout �U  0f��U  �g��U  �iSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �t��U  S�k[.�  ��}&/       Workout     0���U  ����U  0�justforfun_justforfun_ ��U  ����U  0���U  ���U  ����U  Qx�[.�  R�}&/       Birthday    @\��U   ]��U  �]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �b��U  T�	\.�  6�}&/      Workout �U  0f��U  �g��U  �ijustforfun_justforfun_ ��U  �p��U  �q��U  �s��U  �t��U  䍋\.�  p~&/      Workout     л��U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  �W].�  �<~&/       Meeting     p���U  0���U  ��justforfun_justforfun_ _ �U  0���U  ���U  ����U  p���U  �*].�  @~&/      Some_stuffs p��U  0��U  0Some_stuffs_Some_stuffs_ �U   +��U  �+��U  �/��U  p0��U  ,b�].�  mc~&/      Birthday U  ����U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  &��].�  �c~&/       Some_stuffs E��U  �E��U  PFSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �J��U  �].�   e~&/       Appointment p���U  ���U  ��This_stuffs_This_stuffs_ �U  ���U  ����U  @���U  ����U  �+�].�  i~&/       Workout �U  pR��U  �R��U  �SThis_stuffs_This_stuffs_ �U  `V��U   W��U  �W��U  �X��U  ���].�  k~&/       Some_stuffs �H��U  @I��U  �ISome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �M��U  Jc�].�  ]k~&/       Birthday    ����U  `���U  ��Some_stuffs_Some_stuffs_ �U  ����U  `���U  е��U  ����U  ��].�  �k~&/       Meeting     @t��U  �t��U  �uThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Pz��U  �h^.�  ��~&/      Workout     ���U  ����U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ���^.�  l�~&/       Appointment p��U  0��U  0Some_stuffs_Some_stuffs_ �U   +��U  �+��U  �/��U  p0��U  +��^.�  )�~&/       Birthday fs Ю��U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  ��^.�  ��~&/       Birthday nt @��U   ��U  �justforfun_justforfun_ _ �U   	��U  �	��U  @
��U  �
��U   �^.�  Է~&/       Some_stuffs �%��U  0&��U  �&justforfun_justforfun_ ��U  �)��U  0*��U  �*��U  p+��U  	>�.�  ���&/       Appointment p���U  0���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U   .K�.�  ��&/       Meeting     ���U  ���U  0justforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U  @��U  8��.�  �&/       Appointment p���U  0���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p��U  ��t�.�  D؉&/       Some_stuffs ���U  p��U  0justforfun_justforfun_ _ �U  0��U  ���U  0��U  ���U  {�.�  �ى&/       Workout     `\��U  �\��U  �]Some_stuffs_Some_stuffs_ �U  �_��U  p`��U  �`��U  �a��U  �r|�.�  :ډ&/       Some_stuffs е��U  ����U  �This_stuffs_This_stuffs_ �U  ����U  ����U  ���U  ����U  ��.�  ۉ&/       Some_stuffs P���U  ���U  ��This_stuffs_This_stuffs_ �U  p���U  0���U  ����U  0���U  ���.�  lۉ&/       Birthday U  ��	��U   �	��U  ��	This_stuffs_This_stuffs_ �U  ��	��U  P�	��U  ��	��U  P�	��U  :���.�  �݉&/       Meeting ent P���U  ���U  ��justforfun_justforfun_ ��U  ����U  ����U  P���U  ���U  H0�.�  }��&/       Some_stuffs                    justforfun_justforfun_                                       ���.�  	�&/      Appointment �}��U  ����U  pjustforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U  ���U  H���.�  �)�&/       Birthday     c��U  �c��U  `dSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   i��U  �o��.�  Z*�&/       Workout     `���U  ����U  `�This_stuffs_This_stuffs_ �U  `���U   ���U  ����U  `���U  F-��.�  �*�&/      Some_stuffs  ��U  ���U  �This_stuffs_This_stuffs_ �U  0��U  ���U   $��U  �%��U  IE;�.�  �L�&/       Appointment `y��U   z��U  �zThis_stuffs_This_stuffs_ �U  �}��U  ����U  p��U  0���U  \LC�.�  �N�&/      Some_stuffs                    Some_stuffs_Some_stuffs_                                     �"Q�.�  6R�&/       Appointment �	��U  @	��U  �	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �	��U  �o،.�  �t�&/       Some_stuffs                    This_stuffs_This_stuffs_                                     nc�.�  n��&/      Birthday     ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ж��U  �xt�.�  ˜�&/       Meeting     p���U  ���U  ��This_stuffs_This_stuffs_ �U  0���U  ����U  ����U  0���U  �t�.�  ~Ŋ&/      Meeting     �,��U  �-��U  @.This_stuffs_This_stuffs_ �U   1��U  �1��U  �2��U   3��U  B|��.�  (�&/       Some_stuffs 0���U  ���U  ��justforfun_justforfun_ ��U  ����U  0���U  ���U  p���U  ݜ��.�  ��&/      Some_stuffs pF��U  0G��U  �Gjustforfun_justforfun_ ��U  0J��U  �J��U  �K��U  0L��U  �ñ�.�  �&/       Some_stuffs 0"��U  �<��U  0$Some_stuffs_Some_stuffs_ �U  �&��U  �'��U  0(��U  �(��U  �&2�.�  ��&/       Appointment                    This_stuffs_This_stuffs_                                     �?�.�  n�&/      Meeting �U  P[��U  \��U  �`Some_stuffs_Some_stuffs_ �U   l��U  �l��U  �g��U  �h��U  �bۏ.�  6:�&/       Meeting     ����U  p���U  0�This_stuffs_This_stuffs_ �U  ����U  ����U  ����U   ���U  ��ޏ.�  ;�&/       Some_stuffs ����U  ����U  �This_stuffs_This_stuffs_ �U  ����U  `���U  @���U  ���U  9��.�  S=�&/       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             h�r�.�  �`�&/       Some_stuffs ���U  ����U  �This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  �B~�.�  �c�&/      Workout      E��U  �F��U  0KSome_stuffs_Some_stuffs_ �U  �U��U  �V��U  P[��U  \��U  *���.�  ɂ�&/       Workout     ���U  ����U  P�This_stuffs_This_stuffs_ �U  P���U  ����U  P���U  ���U  ���.�  g��&/      Meeting     @]��U   ^��U  �^Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �b��U   ��.�  ���&/       Some_stuffs �p��U   q��U  �wSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �v��U  ɳ��.�  ���&/       Meeting     ���U  `��U  justforfun_justforfun_ ��U   ��U  ���U  ���U  ���U  �Y��.�  �&/       Meeting  nt ��	��U  �	��U  ��	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �	��U  _��.�  9��&/      Workout     0~��U  �~��U  `yThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��@�.�  G׋&/      Meeting ffs ���U  0��U  �Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ���U  �4ǒ.�  ���&/      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             1ns�.�  �%�&/       Workout     ����U  0���U  P
This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  �kx�.�  '�&/       Some_stuffs �w��U  �x��U  PsSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �~��U  (=��.�  It�&/       Appointment `o��U   p��U  �pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �u��U  ��!�.�  㓌&/       Meeting �U  �t��U  �u��U  vThis_stuffs_This_stuffs_ �U  `y��U   z��U  �z��U  `{��U  %�"�.�  8��&/      Some_stuffs  o��U  �o��U  �pjustforfun_justforfun_ ��U  Ps��U  t��U  �t��U  �u��U  �'/�.�  V��&/       Appointment �>��U  ?��U  �?justforfun_justforfun_ _ his_stuffs_This_stuffs_ �U  �D��U  )	��.�  ��&/       Meeting ent  ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  L��.�  �&/      Birthday    @N��U  �N��U  pOSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   S��U  ���.�  �1�&/       Some_stuffs �Y��U   Z��U  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @_��U  l���.�  2�&/      Birthday U  Р��U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  "z��.�  �3�&/       Appointment �	��U   	��U  �	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0#	��U  9���.�  �8�&/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��*�.�  �Z�&/      Some_stuffs P���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �-�.�  �[�&/       Birthday    0���U  ���U  p�justforfun_justforfun_ ��U  ���U  @���U  ���U  ����U  �k<�.�  W_�&/       Appointment ����U  P���U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  �TƘ.�  ���&/       Meeting �U  @���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��Ș.�  E��&/       Workout     0���U   ���U  @�justforfun_justforfun_ ��U  p���U  0���U  ����U  `���U  C*Ϙ.�  脍&/       Appointment ����U  ����U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �Ԙ.�  )��&/      Some_stuffs  ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ж��U  ��՘.�  ���&/       Workout ent ����U  @���U  ��Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ����U  ��V�.�  ���&/       Birthday    0���U  ���U  ��justforfun_justforfun_ _ �U  p���U  ���U  ����U  p���U  �\�.�  ���&/       Some_stuffs P���U  Т��U  ��justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U   ���U  �(c�.�  ˪�&/       Some_stuffs @���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  !:f�.�  ���&/       Appointment 0���U  ����U  0�Some_stuffs_Some_stuffs_ �U  ����U  p���U  ���U  @���U  ���.�  �э&/      Workout ffs ����U  0���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  ���.�  �Ӎ&/       Appointment `V��U   W��U  �WSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   ]��U  ʀ�.�  ��&/       Workout     е��U  ����U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �섚.�  ��&/       Birthday    Н��U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �c��.�  ���&/       Appointment p���U  0���U  ��Some_stuffs_Some_stuffs_ �U  @���U   ���U  ����U  ����U  @��.�  ���&/       Meeting     �7��U  `8��U   9justforfun_justforfun_ ��U  �;��U  `<��U  �<��U  �=��U  G,��.�  (��&/       Meeting     �	��U  0
��U  �
justforfun_justforfun_ ��U  ���U  0��U  ���U  ���U  �ᚚ.�  ���&/       Meeting     ���U  p��U  0This_stuffs_This_stuffs_ �U  ���U  0��U  ���U  ���U  aP��.�  ���&/       Workout     ����U  `���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  >���.�  ��&/      Some_stuffs ����U  `���U  ��This_stuffs_This_stuffs_ �U  ����U  `���U  е��U  ����U  ��&�.�  p�&/      Birthday    ����U  @���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  kX��.�  �ɘ&/       Workout     ���U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  y���.�  �͘&/       Appointment Ъ��U  ����U  P�justforfun_justforfun_ ��U  Ю��U  ����U  ���U  ����U  "E��.�  tИ&/       Appointment  c��U  �c��U  `djustforfun_justforfun_ _ �U  �f��U  �g��U  `h��U   i��U  
��.�  �ј&/      Appointment ���U  ����U  0�This_stuffs_This_stuffs_ �U   ���U  ����U  ����U  @���U  Ī��.�  <��&/      Some_stuffs p���U  0���U  ��justforfun_justforfun_ ��U  p��U  ���U  ���U  p��U  d��.�  <�&/       Appointment ���U  ����U  `�Some_stuffs_Some_stuffs_ �U  ����U  @���U  ����U  @���U  *e�.�  I�&/       Meeting     @f��U  �f��U  @gSome_stuffs_Some_stuffs_ �U  �i��U  @j��U   k��U  �k��U  	��.�  u�&/       Birthday    ���U  Ш��U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  ��.�  x�&/       Workout     � ��U  �!��U  p"Some_stuffs_Some_stuffs_ �U  0%��U  �3��U  @'��U   (��U  $�!�.�  8�&/      Some_stuffs                    This_stuffs_This_stuffs_                                     ���.�  �B�&/      Appointment �	��U  ��	��U  �	Some_stuffs_Some_stuffs_ �U  p�	��U  �	��U  p�	��U   �	��U  x\��.�  �E�&/       Workout     ����U  @���U  ��justforfun_justforfun_ ��U   ���U  ����U   ���U  ����U  ��5�.�  �e�&/       Birthday    p���U  0���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  
�:�.�  g�&/       Meeting     ���U  ����U  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �D�.�  ~i�&/      Appointment ����U  `���U  ��Some_stuffs_Some_stuffs_ �U  ���U  `��U  ��U  ���U  ���.�  ��&/      Birthday                       justforfun_justforfun_                                       ��d�.�  T��&/      Appointment �w��U  �x��U  PsSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �~��U  A��.�  h��&/       Meeting     `h��U   i��U  �iThis_stuffs_This_stuffs_ �U  �l��U  `m��U   ��U  ���U  �L��.�  x��&/       Meeting ffs 0���U  ����U  p�justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  ����U  �} �.�  Cۙ&/       Appointment  $��U  �%��U   +This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �:��U  �$	�.�  zݙ&/      Meeting     ����U  p���U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  7�.�  ��&/       Some_stuffs �K��U  0L��U  �LSome_stuffs_Some_stuffs_ �U  �O��U  pP��U  �P��U  �Q��U  "��.�  ��&/       Meeting                        This_stuffs_This_stuffs_                                     9,��.�  S�&/       Workout     ��U  ���U  �Some_stuffs_Some_stuffs_ �U  ���U  ���U  p��U  0��U  2	��.�  ��&/       Meeting     ����U  P���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  4H��.�  �&/      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             -�D�.�  M.�&/      Some_stuffs ���U  0 ��U  � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0&��U  �bL�.�  :0�&/       Appointment е��U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �n��.�  =P�&/      Appointment ����U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  /j�.�  dy�&/      Meeting     ����U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  p���U  0���U  ����U  ��n�.�  �z�&/       Workout                        This_stuffs_This_stuffs_                                     Pv�.�  |�&/       Birthday    0���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  C�z�.�  �}�&/       Some_stuffs ���U  p��U  0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p!��U  rG|�.�  ~�&/       Birthday    ���U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  ����.�  p��&/      Some_stuffs �t��U  �u��U  vjustforfun_justforfun_ ��U  `y��U   z��U  �z��U  `{��U  � 
�.�  N��&/       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             I՗�.�  �ƚ&/       Birthday    Ц��U  ����U  �Some_stuffs_Some_stuffs_ �U  Ъ��U  ����U  P���U  ���U  |Z��.�  �ƚ&/      Birthday    0���U   ���U  @�This_stuffs_This_stuffs_ �U  p���U  0���U  ����U  `���U  ��E�.�  &�&/      Meeting     ����U  ���U  ЮSome_stuffs_Some_stuffs_ �U  P���U  ���U  ����U  ���U  �K�.�  ���&/       Workout     ���U  ����U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  Y;��.�  �&/       Meeting     �R��U  PS��U  Tjustforfun_justforfun_ ��U  �q��U  `r��U   W��U  �W��U  *l��.�  ��&/       Meeting     ����U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  0���.�  ^�&/       Some_stuffs @b��U  �b��U  �cSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �g��U  h�j�.�  1>�&/       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             YEk�.�  G>�&/       Meeting     P���U  ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  ���.�  �d�&/       Workout     �%��U  0&��U  �&This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p+��U  ��.�  �f�&/       Workout     ����U  p���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  �S�.�  h�&/      Workout     ����U  P���U  �Some_stuffs_Some_stuffs_ �U  P���U  ����U  ����U  P���U  ����.�  ���&/      Some_stuffs �l��U  `m��U   Some_stuffs_Some_stuffs_ �U  �p��U  �q��U  0r��U  �r��U  Yr��.�  g��&/       Workout     `5��U  �5��U  `6This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ;��U  z��.�  ۍ�&/       Birthday    �4��U  p5��U  �9This_stuffs_This_stuffs_ �U   E��U  �F��U  0K��U  �K��U  �6�.�  ٳ�&/      Appointment ����U  ����U  НThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  0���U  ����.�  0֛&/       Some_stuffs 0���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ,���.�  �ܛ&/      Workout     л��U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  1�V�.�  ���&/       Meeting     �+��U   ,��U  �,Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �1��U  �X[�.�  ���&/       Appointment �i��U  pj��U  0kThis_stuffs_This_stuffs_ �U  pm��U  0n��U  �n��U  po��U  
Qu�.�  u�&/       Some_stuffs `���U  ����U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �x�.�  '�&/      Workout     ����U  `���U   �This_stuffs_This_stuffs_ �U  Т��U  P���U  ���U  ����U  p��.�  f%�&/       Meeting                        justforfun_justforfun_                                       ]���.�  �%�&/      Some_stuffs �.��U  @/��U  �/Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �3��U  Z���.�  G&�&/       Birthday    ���U  ����U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  �O��.�  �'�&/       Appointment �{��U  0|��U  �|justforfun_justforfun_ ��U  `���U  ����U  `���U   ���U  ��.�  �O�&/      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �2 �.�  �r�&/      Some_stuffs ���U  ����U  P�This_stuffs_This_stuffs_ �U  P���U  ����U  P���U  ���U  x�/�.�  �v�&/       Appointment @
��U  �
��U  @Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  @��U  ����.�  h��&/      Appointment ����U  P���U  �justforfun_justforfun_ ��U  ���U  p���U  ����U  ����U  `��.�  \��&/       Birthday    �
��U  ���U  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0��U  ����.�  .��&/       Meeting     0���U  ���U  ��justforfun_justforfun_ ��U  p���U  0���U  ����U  0���U  [���.�  ���&/       Birthday nt pG��U  �G��U  �HSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  pL��U  �9X�.�  �&/      Birthday                       justforfun_justforfun_ _Some_stuffs_Some_stuffs_             qij�.�  Fǜ&/       Birthday U   ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  Y���.�  ��&/       Some_stuffs �*��U  p+��U  0,Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �0��U  ���.�  �&/       Appointment  	��U  �	��U  P	justforfun_justforfun_ 	��U  �	��U   	��U  �	��U    	��U  �d��.�  ��&/       Birthday    ����U  @���U  ��Some_stuffs_Some_stuffs_ �U  0���U  ����U  0���U  ����U  <�.�  W�&/      Appointment ���U  p��U  0Some_stuffs_Some_stuffs_ �U  ���U  0 ��U  � ��U  �!��U  �V��.�  �&/       Meeting     ���U  0 ��U  � justforfun_justforfun_ _ �U  �#��U  p$��U  0%��U  �3��U  �՗�.�  p�&/      Meeting     ���U  p��U  0This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �!��U  Q��.�  ��&/       Some_stuffs  |��U  �|��U  �}This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0���U  S;/�.�  2;�&/       Some_stuffs �7	��U   8	��U  �8	This_stuffs_This_stuffs_ �U  �:	��U  `;	��U  <	��U  �<	��U  ��1�.�  �;�&/      Appointment p��U  0��U  0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p0��U  ��2�.�  <�&/       Some_stuffs ��U  ���U  �justforfun_justforfun_ ��U  ���U  ���U  p��U  0��U  ��6�.�  =�&/       Workout     �%��U  0&��U  �&Some_stuffs_Some_stuffs_ �U  �)��U  0*��U  �*��U  p+��U  b�t /�  |�&/       Some_stuffs ����U  p���U  0�justforfun_justforfun_ ��U  ����U  p���U  ����U  ����U  \�t /�  ��&/      Birthday     ���U  ����U  ��justforfun_justforfun_ ��U  ����U  `���U   ���U  ����U  ��w /�  E�&/       Meeting     ����U  p���U  0�This_stuffs_This_stuffs_ �U  ����U  0���U  ���U  ����U  �/�  G5�&/      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             R�/�  r6�&/       Appointment �c��U  @d��U  �dSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   i��U  A�'/�  H;�&/       Birthday nt �2��U   3��U   4This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  `8��U  �̜/�  KY�&/       Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             }�/�  _�&/      Some_stuffs  ��U  ���U  `justforfun_justforfun_ _ �U  `��U   ��U  ���U   ��U  �9/�  n��&/      Meeting      ���U  ����U  `�This_stuffs_This_stuffs_ �U  ����U  `���U  `���U   ���U  alI/�  |��&/       Workout     ����U  `���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U   ��/�  ԧ�&/       Workout �U  �|��U  �}��U  0~This_stuffs_This_stuffs_ �U  `���U   ���U  ����U  `���U  ���/�  %��&/       Appointment @���U   ���U  ��justforfun_justforfun_ ��U  ����U  @���U   ���U  ����U  ���/�  s��&/      Workout     ���U  `��U  justforfun_justforfun_ ��U   ��U  ���U  ���U  ���U  �a�/�  ���&/       Appointment p��U  ���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p$��U  �q/�  )Ѩ&/      Workout     ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  �/�  ���&/       Workout     �<��U  �=��U   >justforfun_justforfun_ ��U  �N��U  PO��U  0A��U  �A��U  O�/�  !��&/      Birthday    ���U  ����U  0�Some_stuffs_Some_stuffs_ �U   ���U  ����U  ����U  @���U  �/�  `��&/       Workout                        This_stuffs_This_stuffs_                                     ��!/�  l��&/       Appointment 0f��U  �g��U  �iThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �t��U  h�/�  ��&/       Appointment ���U  p��U  0This_stuffs_This_stuffs_ �U  ���U  0 ��U  � ��U  �!��U  q��/�  ��&/       Workout     ����U  @���U  ЋThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  6a�/�  �!�&/      Some_stuffs p��U  0��U  0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p0��U  ��/�  �$�&/       Workout     0���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  ��D/�  �H�&/      Birthday    ���U   ��U  �This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  ���U  $y�/�  �n�&/      Appointment ���U  ����U  P�justforfun_justforfun_ ��U  ���U  ����U  ����U  P���U  ��b/�  +��&/       Workout     �e��U  `f��U  �fThis_stuffs_This_stuffs_ �U  �i��U  �j��U  `k��U   l��U  A'n/�  ��&/       Some_stuffs 0A��U  �A��U  �BSome_stuffs_Some_stuffs_ �U  0E��U  �E��U  pF��U  0G��U  K1z/�  ��&/       Appointment 00��U  �0��U  p1This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �5��U  �p�/�  {��&/      Workout                        Some_stuffs_Some_stuffs_                                     -��/�  ���&/      Workout     `/	��U  �/	��U  `0	Some_stuffs_Some_stuffs_ �U  `2	��U  �2	��U  `3	��U  �3	��U  p /�  ���&/       Some_stuffs ����U  @���U  �justforfun_justforfun_ ��U  P���U  ���U   ���U  ����U  �=�/�  �&/       Workout     ���U  0 ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �3��U  �Z�/�  ��&/       Meeting �U  � ��U  �!��U  p"justforfun_justforfun_ ��U  0%��U  �3��U  @'��U   (��U  
�/�  5�&/       Meeting �U  ����U  0���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  { �/�  {�&/       Meeting     �i��U  pj��U  0kSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  po��U  �C�/�  �/�&/      Some_stuffs ����U  `���U   �Some_stuffs_Some_stuffs_ �U  ����U  p���U  0���U  ����U  1��/�  �1�&/       Workout ent ���U  ����U  ��This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  ����U  `zp	/�  <Z�&/       Appointment ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  5nv	/�  �[�&/      Some_stuffs @���U   ���U  ��Some_stuffs_Some_stuffs_ �U  ����U  @���U   ���U  ����U  �a�	/�  B|�&/       Meeting     p:��U  0;��U  �;Some_stuffs_Some_stuffs_ �U  �=��U  �>��U  p?��U  �?��U  @O�	/�  ~�&/       Workout                        justforfun_justforfun_                                       =�	/�  7~�&/      Meeting                        justforfun_justforfun_                                       
/�  8��&/       Some_stuffs ����U  ���U  ЮSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ��
/�  L��&/       Appointment ����U  ����U  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  �9�
/�  �&/      Appointment ���U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ���
/�  ���&/       Birthday    ����U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  `ܭ
/�  |��&/       Appointment p��U  0��U  0justforfun_justforfun_ _ �U   +��U  �+��U  �/��U  p0��U  �,/�  �˪&/       Meeting ffs �R��U   S��U  �SSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  X��U  �;/�  �Ϫ&/      Appointment �&��U  �'��U  0(This_stuffs_This_stuffs_ �U  �*��U  p+��U  0,��U  �,��U  y�D/�  Ҫ&/       Some_stuffs w��U  �w��U  xSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �|��U  $Z�/�  ���&/      Meeting     0��U  ���U  �This_stuffs_This_stuffs_ �U  ���U  p��U  0��U  ���U  x�n/�  [�&/       Appointment ����U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P��U  �+q/�  �&/      Workout      ���U  ����U  0�justforfun_justforfun_ _ �U  ����U  P���U  ����U  P���U  ��x/�  � �&/       Some_stuffs ���U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0���U  0{�/�  �?�&/       Meeting     е��U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  y,/�  �G�&/       Meeting     � ��U  �!��U  p"justforfun_justforfun_ ��U  0%��U  �3��U  @'��U   (��U  ���/�  6i�&/       Appointment v��U  �v��U  0~This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �|��U  ��/�  �i�&/       Meeting     pm��U  0n��U  �nThis_stuffs_This_stuffs_ �U  pq��U  �q��U  pr��U  �r��U  ��/�  nj�&/      Some_stuffs  E��U  �F��U  0KSome_stuffs_Some_stuffs_ �U  �U��U  �V��U  P[��U  \��U  !/�  ���&/       Birthday    p?��U  �?��U  p@This_stuffs_This_stuffs_ �U  pB��U  �B��U  �C��U  0D��U  \�#/�  K��&/      Birthday U   o��U  �o��U  �pSome_stuffs_Some_stuffs_ �U  Ps��U  t��U  �t��U  �u��U  ˠ-/�  ͐�&/       Meeting     �		��U  `
	��U  �
	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �	��U  ��0/�  ���&/       Birthday     ���U  ����U  ��justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  p���U  �$�/�  ̵�&/       Birthday    ����U  ����U  p�This_stuffs_This_stuffs_ �U  ����U  @���U  ����U  ����U  ��/�  ���&/       Appointment ����U  `���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  ��/�  P��&/      Workout     ����U  ����U  @�Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  @���U  ��/�  ּ�&/       Workout     ����U  0���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �r�/�  ���&/       Birthday     4��U  �4��U  `5This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �9��U  ��h/�  ��&/       Meeting     ����U  P���U  �This_stuffs_This_stuffs_ �U  `���U   ���U  ���U  ����U  \�s/�  K�&/      Some_stuffs                    justforfun_justforfun_                                       u/�  ��&/       Meeting �U  0f��U  �g��U  �iSome_stuffs_Some_stuffs_ �U  �p��U  �q��U  �s��U  �t��U  �M�/�  n�&/       Birthday    0���U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  l��/�  ��&/      Appointment ����U  @���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  Ae�/�  ��&/       Birthday    ����U  ����U  ��justforfun_justforfun_ ��U  ����U  @���U   ���U  ����U  �/�  �	�&/       Meeting     p��U  0��U  �This_stuffs_This_stuffs_ �U  �	��U  0
��U  �
��U  ���U  xf�/�  ;0�&/       Birthday     ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  a"%/�  <S�&/       Workout      ���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  `���U  ����U  `���U  ��1/�  oV�&/      Appointment ����U  P���U  �Some_stuffs_Some_stuffs_ �U  `���U   ���U  ���U  ����U  