>~
 /   d~
 /      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ݦ
 /   ��
 /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ��
 /   ��
 /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     $ /   [ /      Birthday     ��/V  @��/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  C /   6C /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     � /   �� /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               �� /   �� /      Birthday    �		�/V  �
	�/V  	Some_stuffs_Some_stuffs_ /V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  5� /   �� /      Some_stuffs  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  � /   n /      Meeting /V  p��/V  ���/V  ��This_stuffs_This_stuffs_ /V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  2) /   _) /      Meeting &V  �(Կ&V  P*Կ&V  �/�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   ;Կ&V  �<Կ&V   EԿ&V  �@Կ&V   BԿ&V  @CԿ&V  �JԿ&V  `FԿ&V  �GԿ&V  `IԿ&V  �PԿ&V   LԿ&V  @MԿ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  {O /   �S /       Appointment PIӿ&V  �Jӿ&V  �M�Some_stuffs_Some_stuffs_ &V  �Vӿ&V  @Xӿ&V  p[ӿ&V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  9{ /   H{ /      Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  6� /   g� /       Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �� /   �� /      Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  B /    /      Workout     ���/V  ���/V   �This_stuffs_This_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  �= /   �= /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �� /   �� /   	   Appointment ���/V   ��/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �/V  P�/V  ��/V  �/V  ɱ /   /� /   	   Some_stuffs  ��/V  @��/V  ��Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  �� /   �� /      Meeting     ���/V  ���/V  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  7� /   $� /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �* /   p' /      Birthday V  � �/V  0�/V  pjustforfun_justforfun_ �/V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  �Q /   R /      Workout     �!�/V  #�/V  �Some_stuffs_Some_stuffs_ /V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V  0q /   3p /      Appointment P$�/V  �%�/V   'justforfun_justforfun_ �/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  �� /   �� /       Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               �� /   �� /      Appointment �/�/V   1�/V  �5Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  P��/V  ���/V  `��/V   ��/V  Q� /   V� /      Meeting /V  �
�/V  

�/V  �
justforfun_justforfun_ 
�/V   
�/V  `
�/V  �
�/V  
�/V  P
�/V  �
�/V  P
�/V  �
�/V  �
�/V  
�/V  P
�/V  � 
�/V  "
�/V  :
�/V   '
�/V  `(
�/V  �)
�/V  �*
�/V   ,
�/V  �-
�/V   /
�/V  `0
�/V  �1
�/V  `3
�/V  �4
�/V   6
�/V  �7
�/V  �N
�/V  P;
�/V  �[ /   �[ /   	   Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �~ /   �~ /      Appointment ���/V   ��/V  `�Some_stuffs_Some_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  Х /   � /      Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             � /   '� /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             5� /   :� /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ~ /   � /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �o /   �o /      Meeting     �R�/V  �S�/V  UThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  �� /   �� /      Appointment  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  f� /   �� /      Appointment ���/V   ��/V  ��Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  � /   � /      Birthday    ���/V   ��/V  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  �1 /   �. /      Appointment �	�/V  0�	�/V  p�	Some_stuffs_Some_stuffs_ /V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  p�	�/V  @�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  �W /   �W /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �� /   ¤ /      Some_stuffs ��/V  `�/V  �#Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  � /   '� /      Meeting     `��/V  ���/V  0�This_stuffs_This_stuffs_ /V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  k� /   � /      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ! /   A /      Appointment p��/V  ��/V  0�justforfun_justforfun_ �/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  p�/V  p�/V  |D /   �D /      Appointment ���/V  Ъ�/V  P�justforfun_justforfun_ �/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V  Q� /   h� /      Birthday V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V   /   E /      Appointment @��/V  ���/V  ��This_stuffs_This_stuffs_ /V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  r' /   �' /      Meeting &V  ��ӿ&V  P�ӿ&V  ���This_stuffs_This_stuffs_ &V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  ��( /   ��( /      Meeting     `��/V  ��/V  `�justforfun_justforfun_ �/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  `��/V  0��/V  p��/V  ���/V   ��/V  `��/V  ���/V  0��/V  �%) /   �') /       Birthday    �#�/V  P%�/V  �)This_stuffs_This_stuffs_ /V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  �t) /   �t) /      Workout     ���/V  ���/V  �Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  Н) /   ��) /      Birthday V  PZ	�/V  �[	�/V  `L	This_stuffs_This_stuffs_ /V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  E�) /   J�) /      Meeting     �	�/V  �/V  Pjustforfun_justforfun_ �/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �* /   �* /      Some_stuffs ���/V  ���/V   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  �5* /   �5* /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �* /   q�* /       Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               ��* /   Ы* /      Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ��* /   ��* /      Some_stuffs `M�/V  �N�/V  �ZSome_stuffs_Some_stuffs_ /V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  K+ /   ��* /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �"+ /   a#+ /      Meeting /V  �z�/V  ���/V  �~Some_stuffs_Some_stuffs_ /V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  aH+ /   wH+ /   	   Some_stuffs Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  �r+ /   s+ /      Workout /V   <�/V  �F�/V  @?This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  ��+ /   )�+ /   	   Birthday    ��/V   �/V  �!justforfun_justforfun_ �/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  ��+ /   "�+ /   	   Meeting /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  _�+ /   v�+ /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �[, /   (^, /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �, /   �, /   	   Meeting     ���/V  ���/V   �justforfun_justforfun_ �/V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  ��, /   ��, /       Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �, /   9�, /       Meeting     P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �B- /   �G- /      Meeting     P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �r- /   �r- /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               �?8 /   �?8 /      Some_stuffs ���/V  @��/V  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  �f8 /   0g8 /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��8 /   ��8 /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               $9 /   l9 /      Appointment ���/V  P��/V  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V  h-9 /   p-9 /   	   Birthday    P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  !R9 /   �W9 /      Meeting     `	�/V  �	�/V  	This_stuffs_This_stuffs_ /V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  ţ9 /   ��9 /       Some_stuffs ���/V   ��/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  ��9 /   ��9 /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �: /   �: /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �c: /   �f: /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ��: /   ܏: /   	   Some_stuffs �W�/V  �X�/V  �eThis_stuffs_This_stuffs_ /V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V   �: /   '�: /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     -+; /   �(; /      Appointment p`
�/V  �a
�/V  �z
justforfun_justforfun_ 
�/V  i
�/V  Pj
�/V  �k
�/V  �l
�/V  n
�/V  Po
�/V  �p
�/V  Pr
�/V  �s
�/V  u
�/V  �v
�/V  �w
�/V  y
�/V  �
�/V  0}
�/V  p~
�/V  �
�/V  ��
�/V  0�
�/V  p�
�/V  ��
�/V  ��
�/V  0�
�/V  ��
�/V  ��
�/V   �
�/V  ��
�/V   �
�/V  `�
�/V  \U; /   �U; /      Workout /V  �	�/V  P�	�/V  ��	This_stuffs_This_stuffs_ /V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  Ю	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  fu; /   �u; /      Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               ^�; /   w�; /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               $�; /   ��; /      Some_stuffs �
�/V  
�/V  P
Some_stuffs_Some_stuffs_ /V   '
�/V  `(
�/V  �)
�/V  �*
�/V   ,
�/V  �-
�/V   /
�/V  `0
�/V  �1
�/V  `3
�/V  �4
�/V   6
�/V  �7
�/V  �N
�/V  P;
�/V  �<
�/V  >
�/V  �?
�/V  A
�/V  PB
�/V  �C
�/V  �D
�/V  F
�/V  PG
�/V  �H
�/V  �I
�/V  K
�/V  �L
�/V  �c
�/V  ]�; /   ��; /      Workout     P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  +< /   �< /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ;< /   A;< /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �^< /   �^< /      Birthday V   �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  -�< /   P�< /      Appointment ���/V  Д�/V  �This_stuffs_This_stuffs_ /V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  h�< /   ��< /      Appointment ��	�/V  Щ	�/V  �	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  XaG /   �aG /      Birthday V  `	�/V  �	�/V  	This_stuffs_This_stuffs_ /V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  ԨG /   �G /      Birthday    ���/V  0��/V  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  �G /   ��G /      Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  iH /   �H /      Appointment ���/V   ��/V  `�This_stuffs_This_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  ��H /   ��H /      Workout     PIӿ&V  �Jӿ&V  �M�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �H /   <�H /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �2I /   �2I /      Appointment ��/V  `�/V  �#This_stuffs_This_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  _I /   YI /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     p�I /   ��I /      Birthday    ���/V  ���/V   �This_stuffs_This_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  :�I /   :�I /      Appointment ��Կ&V   �Կ&V  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  ��Կ&V  `�Կ&V  ��Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  `�Կ&V  0�Կ&V  p�Կ&V   �Կ&V  @�Կ&V  ��Կ&V   �Կ&V  P�Կ&V  ��Կ&V  �Կ&V  0�Կ&V  p�Կ&V  �Կ&V  `�Կ&V  ��Կ&V  ЩԿ&V  �Կ&V  P�Կ&V  ��Կ&V  �Կ&V  �I /   ��I /      Appointment ��	�/V  ��	�/V   �	Some_stuffs_Some_stuffs_ /V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  	"J /   �J /       Appointment @	�/V  �,	�/V  �	Some_stuffs_Some_stuffs_ /V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  "iJ /   LiJ /      Birthday V  ��ӿ&V  p�ӿ&V  0��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  ��J /   ��J /   	   Meeting /V  ���/V  ���/V   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  (�J /   <�J /      Appointment  ��/V  ���/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �SK /   �TK /       Appointment  U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ؠK /   ڠK /      Birthday    �u	�/V  �v	�/V  `x	Some_stuffs_Some_stuffs_ /V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  $�K /   ��K /      Meeting     0H�/V  pI�/V  �JSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  Q�K /   _�K /      Some_stuffs � �/V  0�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  L�V /   l�V /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               p�V /   ��V /      Appointment @B�/V  �C�/V  PSome_stuffs_Some_stuffs_ /V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  6�V /   G�V /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             RW /   �W /      Meeting      <�/V  �F�/V  @?Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  >@W /   N@W /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     paW /   �aW /      Workout     �!�/V  #�/V  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V  ͌W /   όW /       Meeting     ��/V  `�/V  �#Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  O�W /   ɯW /       Workout     �	�/V  �/V  PSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  P�W /   �W /      Meeting     �u	�/V  �v	�/V  `x	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��	�/V   �	�/V  @�	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  � X /   �X /      Appointment `��/V  ���/V  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  �&X /   �&X /      Birthday V  U�/V  PV�/V  �WSome_stuffs_Some_stuffs_ /V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  aMX /   `MX /      Meeting /V  �Z�/V  �[�/V  �RSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V  ��X /   \�X /      Some_stuffs ��/V  P��/V  ��justforfun_justforfun_ �/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ��X /   ��X /      Meeting     PZ	�/V  �[	�/V  `L	Some_stuffs_Some_stuffs_ /V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �X /   ��X /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             {Y /   �Y /      Workout     �#�/V  P%�/V  �)This_stuffs_This_stuffs_ /V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  �<Y /   �<Y /   	   Appointment ���/V   ��/V  `�Some_stuffs_Some_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  q�Y /   (�Y /      Birthday    P�/V  ��/V  This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  ��Y /   `�Y /      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     &Z /   �'Z /      Appointment `FԿ&V  �GԿ&V  `I�This_stuffs_This_stuffs_ &V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  @      �HZ /   cGZ /      Appointment ���/V  ���/V  p�This_stuffs_This_stuffs_ /V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  mqZ /   uqZ /      Meeting /V  ���/V   ��/V  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  G�Z /   ��Z /       Birthday V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  ��Z /   ��Z /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �[ /   �	[ /   	   Some_stuffs ��/V  p�/V  pThis_stuffs_This_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  �
f /   �	f /      Some_stuffs  U�/V  pW�/V  0Yjustforfun_justforfun_ �/V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �.f /   Q1f /      Some_stuffs �z�/V  ���/V  �~Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  }f /   >}f /      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     E�f /   ȣf /      Appointment @��/V  � 	�/V  �	justforfun_justforfun_ 	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  S�f /   >�f /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               =�f /   \�f /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               Xg /   �g /   	   Some_stuffs �		�/V  �
	�/V  	This_stuffs_This_stuffs_ /V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  HBg /   {Bg /      Birthday V  T	�/V  PU	�/V  �V	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  {lg /   Hhg /       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ��g /   2�g /      Some_stuffs P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��g /   ��g /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               ��g /   ��g /      Meeting      ��/V  @��/V  ��This_stuffs_This_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  h /   h /      Meeting /V  `	�/V  �	�/V  	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  �0h /   1h /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �{h /   &xh /      Meeting     P|	�/V  �}	�/V  �m	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  ��h /   �h /      Appointment @3	�/V  �4	�/V  �5	Some_stuffs_Some_stuffs_ /V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  O�h /   ��h /      Meeting     PIӿ&V  �Jӿ&V  �M�Some_stuffs_Some_stuffs_ &V  �Vӿ&V  @Xӿ&V  p[ӿ&V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �h /   ��h /      Meeting     P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �;i /   �;i /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             gi /   gi /      Appointment  ��/V  ���/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  ��i /   ��i /      Meeting     Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  t�i /   ~�i /      Appointment ���/V  Д�/V  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ��i /   �i /      Some_stuffs ���/V  Д�/V  �justforfun_justforfun_ �/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  QPj /   gPj /      Birthday    ��/V  `�/V  �#justforfun_justforfun_ �/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  �uj /   �uj /       Workout &V   �ҿ&V  p�ҿ&V  0��justforfun_justforfun_ ҿ&V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  UPu /   �Pu /      Appointment  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  1ou /   �pu /      Meeting     p��/V  ��/V  0�Some_stuffs_Some_stuffs_ /V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  p�/V  p�/V  ��u /   ��u /      Some_stuffs �z�/V  ���/V  �~This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  ��u /   ��u /       Some_stuffs ���/V  Д�/V  �justforfun_justforfun_ �/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  V�u /   �u /      Some_stuffs P�/V  ��/V  This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �v /   �v /      Workout      ��/V  ���/V  ��This_stuffs_This_stuffs_ /V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �5v /   �5v /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     _v /   1_v /      Appointment `	�/V  �	�/V  	Some_stuffs_Some_stuffs_ /V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  $�v /   K�v /      Workout /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  4�v /   X�v /      Appointment ���/V   ��/V  @�This_stuffs_This_stuffs_ /V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  G�v /   ��v /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             w /   "w /      Birthday    � �/V  0�/V  pjustforfun_justforfun_ �/V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  Ew /   �Hw /      Meeting     ���/V  @��/V  p�Some_stuffs_Some_stuffs_ /V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  �ow /   -mw /       Some_stuffs ��/V  p�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  ��w /   ��w /      Appointment PIӿ&V  �Jӿ&V  �M�This_stuffs_This_stuffs_ &V  �Vӿ&V  @Xӿ&V  p[ӿ&V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �w /   ��w /      Appointment P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  :�w /   X�w /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �x /   Bx /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     \^x /   �^x /      Birthday V  �	�/V  0�	�/V  p�	This_stuffs_This_stuffs_ /V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  p�	�/V  @�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V   �	�/V  `�	�/V  ��	�/V  P�	�/V  ��	�/V  0�	�/V  p�	�/V  9}x /   :}x /      Meeting     �	�/V  �/V  PThis_stuffs_This_stuffs_ /V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  ��x /   �x /      Birthday    ���/V  @��/V  p�This_stuffs_This_stuffs_ /V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  ��x /   �x /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               �y /   �y /      Some_stuffs ���/V   ��/V  `�justforfun_justforfun_ �/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  �ky /   �ky /       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �y /   (�y /      Workout /V  ���/V  ���/V   �justforfun_justforfun_ �/V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  d� /   Fd� /      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ��� /   ʷ� /      Meeting /V  �W�/V  �X�/V  �eSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  �� /   � /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               >z� /   �z� /       Some_stuffs ���/V  @��/V  p�Some_stuffs_Some_stuffs_ /V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  6�� /   5�� /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             w� /   6� /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               }?� /   ~?� /      Meeting /V  ��/V   �/V  �!justforfun_justforfun_ �/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  Ab� /   ub� /      Meeting     ���/V  0��/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  �� /   �� /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     9؆ /   V؆ /      Appointment Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  ��� /   ��� /   	   Appointment  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  s+� /   �"� /       Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �P� /   _J� /      Birthday    PZ	�/V  �[	�/V  `L	Some_stuffs_Some_stuffs_ /V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  ex� /   #q� /      Birthday V  � �/V  0�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  �� /   >�� /      Birthday    �	�/V  �/V  PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �� /   �� /   	   Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     � /   6� /      Workout     ��/V  `�/V  �#justforfun_justforfun_ �/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  �;� /   �;� /      Appointment �#�/V  P%�/V  �)Some_stuffs_Some_stuffs_ /V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  �_� /   �_� /       Appointment p[ӿ&V  �\ӿ&V  0`�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  �� /   m�� /   	   Birthday    �ӿ&V  `�ӿ&V  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  �؈ /   �؈ /   	   Meeting     ���/V   ��/V  `�This_stuffs_This_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  D�� /   ^�� /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �Г /   qՓ /      Appointment P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  Q� /   }� /       Some_stuffs P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �E� /   �E� /      Some_stuffs T	�/V  PU	�/V  �V	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  �m� /   �i� /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               ٓ� /   ٓ� /       Some_stuffs  ��/V  @��/V  ��This_stuffs_This_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  `� /   n� /      Workout     @��/V  � 	�/V  �	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  �-� /   �-� /      Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��� /   ã� /   	   Birthday V  PZ	�/V  �[	�/V  `L	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �˕ /   *̕ /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �� /   �� /      Meeting      ��/V  @��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  �A� /   B� /      Workout     �#�/V  P%�/V  �)Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  �m� /   �m� /      Workout     ��/V  `�/V  �#This_stuffs_This_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  Ҳ� /   㲖 /      Meeting &V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �� /   � /   	   Appointment PIӿ&V  �Jӿ&V  �M�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �W� /   Q� /      Birthday    ���/V  Ъ�/V  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V  T~� /   W~� /       Appointment ��	�/V  ��	�/V   �	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  桗 /   裗 /      Appointment �~�/V   ��/V  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  lŗ /   �ŗ /      Birthday    ���/V  P��/V  �This_stuffs_This_stuffs_ /V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V  �� /   �� /       Some_stuffs ���/V   ��/V  ��Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  �� /   �� /      Workout &V  `FԿ&V  �GԿ&V  `I�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  [=� /   :;� /      Birthday V  0~Կ&V  pԿ&V  �x�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  `�Կ&V  ��Կ&V  @�Կ&V  @�Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  `�Կ&V  0�Կ&V  p�Կ&V   �Կ&V  @�Կ&V  ��Կ&V   �Կ&V  P�Կ&V  ��Կ&V  �Կ&V  0�Կ&V  p�Կ&V  �Կ&V  `�Կ&V  �� /   �� /      Appointment ��/V  `�/V  �#This_stuffs_This_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  &>� /   8>� /      Some_stuffs �ӿ&V  p�ӿ&V  p��This_stuffs_This_stuffs_ &V  �ӿ&V  `�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  �a� /   �a� /      Some_stuffs ���/V  ���/V  �Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  `�� /   :�� /      Meeting     �		�/V  �
	�/V  	justforfun_justforfun_ 	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  � /   �� /      Birthday    �	�/V  �/V  Pjustforfun_justforfun_ �/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  Eף /   wף /      Workout     �	�/V  �/V  PSome_stuffs_Some_stuffs_ /V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  5�� /   �� /      Some_stuffs "
�/V  :
�/V   '
Some_stuffs_Some_stuffs_ /V   ,
�/V  �-
�/V   /
�/V  `0
�/V  �1
�/V  `3
�/V  �4
�/V   6
�/V  �7
�/V  �N
�/V  P;
�/V  �<
�/V  >
�/V  �?
�/V  A
�/V  PB
�/V  �C
�/V  �D
�/V  F
�/V  PG
�/V  �H
�/V  �I
�/V  K
�/V  �L
�/V  �c
�/V  e
�/V  �O
�/V  0Q
�/V  pR
�/V  �(� /   %� /      Meeting     P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  1O� /   :O� /      Appointment  ��/V  @��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  u� /   =o� /      Appointment 0]�/V  p^�/V  �_Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  j�� /   ��� /      Workout &V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  ��� /   N�� /       Some_stuffs  U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �� /   � /      Birthday    ���/V   ��/V  @�This_stuffs_This_stuffs_ /V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   8� /   "8� /      Birthday V  "
�/V  :
�/V   '
This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  `0
�/V  �1
�/V  `3
�/V  �4
�/V   6
�/V  �7
�/V  �N
�/V  P;
�/V  �<
�/V  >
�/V  �?
�/V  A
�/V  PB
�/V  �C
�/V  �D
�/V  F
�/V  PG
�/V  �H
�/V  �I
�/V  K
�/V  �L
�/V  �c
�/V  e
�/V  �O
�/V  0Q
�/V  pR
�/V  ia� /   ha� /      Meeting     ���/V  @��/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  Z�� /   f�� /      Appointment ��ӿ&V  p�ӿ&V  0��This_stuffs_This_stuffs_ &V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  ��� /   ��� /      Birthday    P�/V  ��/V  Some_stuffs_Some_stuffs_ /V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  ]D� /   fD� /      Meeting     ��/V  `�/V  �#justforfun_justforfun_ �/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  �j� /   l� /      Workout     P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  Ք� /   Ք� /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �� /   K� /      Appointment `'	�/V  �(	�/V  �)	This_stuffs_This_stuffs_ /V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  �R	�/V  T	�/V  �Z� /   �Z� /      Appointment �z�/V  ���/V  �~Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  �*� /   �*� /      Birthday V  `M�/V  �N�/V  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  @      �X� /   W� /       Workout     P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  3x� /   �|� /      Some_stuffs PIӿ&V  �Jӿ&V  �M�justforfun_justforfun_ ӿ&V  �Vӿ&V  @Xӿ&V  p[ӿ&V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �� /   P�� /   	   Appointment P�/V  PQ�/V  0HThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  �̲ /   Ͳ /      Workout     0]�/V  p^�/V  �_This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  �� /   ��� /      Some_stuffs ���/V   ��/V  @�This_stuffs_This_stuffs_ /V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  `��/V  0��/V  p��/V  ���/V  0@� /   X@� /       Birthday    �~�/V   ��/V  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  퍳 /   #�� /      Workout     `M�/V  �N�/V  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  K�� /   ݵ� /       Appointment  �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  Tٳ /   0ڳ /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �� /   �� /      Meeting /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  N� /   $N� /      Appointment ��/V  p�/V  pjustforfun_justforfun_ �/V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  �z� /   �z� /       Workout     ��/V  `�/V  �#Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  �� /   �� /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               �Ǵ /   CŴ /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             P� /   z� /      Workout     p�	�/V  ��	�/V  ��	justforfun_justforfun_ 	�/V   �	�/V  `�	�/V  ��	�/V  P�	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  0�	�/V  ��	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  �
�/V  �
�/V  ��	�/V  �	�/V  P 
�/V  �
�/V  
�/V  P
�/V  �
�/V  
�/V  �
�/V  

�/V  �
�/V  E9� /   x9� /       Birthday V  ���/V  P��/V  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V  �^� /   �^� /      Meeting /V   ��/V  `��/V  мThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  X�� /   n�� /      Some_stuffs �	�/V  0�	�/V  p�	Some_stuffs_Some_stuffs_ /V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  p�	�/V  @�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V   �	�/V  `�	�/V  ��	�/V  P�	�/V  ��	�/V  0�	�/V  p�	�/V  J�� /   K�� /      Birthday V  `FԿ&V  �GԿ&V  `I�Some_stuffs_Some_stuffs_ &V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  YԵ /   �Ե /      Birthday    ��	�/V   �	�/V  p�	This_stuffs_This_stuffs_ /V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  p�	�/V  @�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��� /   J�� /   	   Meeting     Ј�/V  P��/V  ЏSome_stuffs_Some_stuffs_ /V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  n$� /   �$� /      Meeting &V  `�Կ&V  ��Կ&V  `��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  p�Կ&V   �Կ&V  @�Կ&V  ��Կ&V   �Կ&V  P�Կ&V  ��Կ&V  �Կ&V  0�Կ&V  p�Կ&V  �Կ&V  `�Կ&V  ��Կ&V  ЩԿ&V  �Կ&V  P�Կ&V  ��Կ&V  �Կ&V  ��Կ&V  �Կ&V  `�Կ&V  ��Կ&V   �Կ&V  ��Կ&V  �Կ&V  �Կ&V  Hu� /   ou� /      Appointment `	�/V  �	�/V  	Some_stuffs_Some_stuffs_ /V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  ��� /   ��� /   	   Workout     ��/V  P��/V  ��This_stuffs_This_stuffs_ /V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ��� /   ��� /      Some_stuffs  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  hrŭ}�  ��
 /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                      ���}�  H{ /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �+�}�  �= /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             0�z�}�  �� /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ��p�}�  �� /       Workout &V  p[ӿ&V  �\ӿ&V  0`�justforfun_justforfun_ ӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  8��}�  �� /      Workout /V  @	�/V  �,	�/V  �	justforfun_justforfun_ 	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V   �A�}�  �[ /   	   Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     X��}�  �~ /      Appointment �ӿ&V  p�ӿ&V  p��Some_stuffs_Some_stuffs_ &V  �ӿ&V  `�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  ����}�  :� /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     P_i�}�  � /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ���}�  ¤ /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     (��}�  Y /      Workout     P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ����}�  h� /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     x�� ~�  E /      Appointment p[ӿ&V  �\ӿ&V  0`�This_stuffs_This_stuffs_ &V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  hd�0~�  �%) /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��{3~�  J�) /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               В_5~�  �5* /      Some_stuffs ��ӿ&V  P�ӿ&V  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  �V7~�  ��* /       Workout     @��/V  ���/V  ��justforfun_justforfun_ �/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V  �~�7~�  ��* /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             XV�9~�  wH+ /   	   Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               ���:~�  s+ /      Workout &V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  8�:A~�  9�, /       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �-�q~�  �?8 /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     Mv~�  /R9 /      Appointment 0s�/V  pt�/V  �uSome_stuffs_Some_stuffs_ /V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  Py�w~�  ��9 /      Meeting     ���/V   ��/V  @�justforfun_justforfun_ �/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  ��{~�  ܏: /   	   Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             Ȍ=~~�  /+; /      Meeting     ��/V  p�/V  pjustforfun_justforfun_ �/V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  �-x�~�  ��; /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��΂~�  A;< /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               ���~�  P�< /      Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ���~�  �H /      Appointment ��ӿ&V  p�ӿ&V  0��This_stuffs_This_stuffs_ &V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  8�ɽ~�  =�I /      Birthday    ��/V  P��/V  ��justforfun_justforfun_ �/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  �ʊ�~�  -"J /      Meeting     �g	�/V  �h	�/V  P|	This_stuffs_This_stuffs_ /V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  ��\�~�  ��J /   	   Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     XQ�~�  _�K /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     H1�~�  όW /       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     0(��~�  �&X /      Birthday V  �ӿ&V  p�ӿ&V  p��Some_stuffs_Some_stuffs_ &V  �ӿ&V  `�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  �xl�~�  `MX /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ��� �  ��Y /      Meeting     Ј�/V  P��/V  ЏSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  8��  uqZ /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �jw:�  \�f /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               `#�<�  ��g /      Some_stuffs P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  (�?>�  ��g /      Meeting     p[ӿ&V  �\ӿ&V  0`�This_stuffs_This_stuffs_ &V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  pղ?�  1h /      Workout &V  �9Կ&V   ;Կ&V  �<�This_stuffs_This_stuffs_ &V  @CԿ&V  �JԿ&V  `FԿ&V  �GԿ&V  `IԿ&V  �PԿ&V   LԿ&V  @MԿ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  �-D�  �;i /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �q�H�  gPj /      Birthday V   �ҿ&V  p�ҿ&V  0��justforfun_justforfun_ ҿ&V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  ��x�  �Pu /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �'�x�  Jou /      Some_stuffs �	�/V  P�	�/V  ��	Some_stuffs_Some_stuffs_ /V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  Ю	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  (�Ky�  ��u /      Some_stuffs p[ӿ&V  �\ӿ&V  0`�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  �3]{�  �v /   	   Appointment �Q	�/V  �R	�/V  T	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  p���  :}x /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �̺��  �ky /       Meeting     �Vӿ&V  @Xӿ&V  p[�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  �S��  (�y /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               ЭE��  ʷ� /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �퇻�  �� /      Some_stuffs �	�/V  P�	�/V  ��	justforfun_justforfun_ 	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  Ю	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V  �����  ~?� /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               �n��  ub� /      Meeting &V   RԿ&V  �SԿ&V   U�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  pԿ&V  �xԿ&V  �yԿ&V  p{Կ&V  �|Կ&V  ��Կ&V   �Կ&V  ��Կ&V  �}*��  �� /      Birthday V   >Կ&V  @?Կ&V  �9�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �JԿ&V  `FԿ&V  �GԿ&V  `IԿ&V  �PԿ&V   LԿ&V  @MԿ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  Ѕi��  V؆ /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               ���  ��� /   	   Appointment ��ӿ&V  p�ӿ&V  0��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  �'n��  �P� /      Appointment ��	�/V  ��	�/V   �	Some_stuffs_Some_stuffs_ /V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  ����  6� /      Workout &V  ��ӿ&V  P�ӿ&V  ���justforfun_justforfun_ ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  H��  �؈ /   	   Meeting &V  �ӿ&V  p�ӿ&V  p��This_stuffs_This_stuffs_ &V  �ӿ&V  `�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  �Wj��  }� /       Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               Hk��  ٓ� /       Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �����  �� /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ��_��  �m� /      Workout &V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  P�e?��  �� /      Birthday V  �9Կ&V   ;Կ&V  �<�justforfun_justforfun_ Կ&V  @CԿ&V  �JԿ&V  `FԿ&V  �GԿ&V  `IԿ&V  �PԿ&V   LԿ&V  @MԿ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  h�@��  wף /      Workout &V   RԿ&V  �SԿ&V   U�Some_stuffs_Some_stuffs_ &V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  pԿ&V  �xԿ&V  �yԿ&V  p{Կ&V  �|Կ&V  ��Կ&V   �Կ&V  ��Կ&V  pc�@��  4�� /      Some_stuffs  U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  PiB��  :O� /      Appointment p[ӿ&V  �\ӿ&V  0`�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  ���F��  ha� /      Meeting &V  PIӿ&V  �Jӿ&V  �M�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  `�mJ��  fD� /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               x�K��  �j� /       Appointment �z�/V  ���/V  �~Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  ؂�K��  Ք� /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �O��  �Z� /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     P��}��  �*� /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     p?���  P�� /   	   Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �H���  Ͳ /      Workout &V  `sԿ&V  �tԿ&V  0~�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   �Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  @�Կ&V  @�Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  `�Կ&V  0�Կ&V  p�Կ&V   �Կ&V  @�Կ&V  ��Կ&V   �Կ&V  P�Կ&V  ��Կ&V  �Կ&V  0�Կ&V  p�Կ&V  X(ۀ��  � /      Meeting     � �/V  0�/V  pThis_stuffs_This_stuffs_ /V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  � ����  ��� /      Appointment ���/V  Д�/V  �justforfun_justforfun_ �/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  0|���  �� /      Meeting &V  ��ӿ&V  P�ӿ&V  ���Some_stuffs_Some_stuffs_ &V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  ������  $N� /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               p����  �z� /       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     P۲���  x9� /       Birthday V  ��ӿ&V  p�ӿ&V  0��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  ��S���  �^� /      Meeting &V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V   M���  �Ե /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ,?���  ��� /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ���,�O d~
 /      Workout     ���/V   ��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  �R�-�O ��
 /      Some_stuffs � �/V  0�/V  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  x+�/�O _) /      Meeting     P$�/V  �%�/V   'This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  ��]0�O g� /       Birthday    ��/V  p�/V  pjustforfun_justforfun_ �/V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  xl�-1�O _ /      Workout     ���/V  ���/V   �Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  �dA3�O "R /      Birthday    �e�/V  �f�/V  0]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  P��H�O � /      Workout     P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �/��I�O �� /   	   Some_stuffs ���/V   ��/V  ��Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �/V  P�/V  ��/V  �/V  (��N�O �' /      Meeting     ���/V   ��/V  `�This_stuffs_This_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  ����d�O Ù+ /      Meeting     ���/V  ���/V  @�justforfun_justforfun_ 	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  h�ѭf�O ��, /       Meeting /V  0s�/V  pt�/V  �uThis_stuffs_This_stuffs_ /V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  ��{�O ��8 /      Meeting     P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  H�.&}�O ��9 /      Meeting /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ���_}�O �: /      Birthday V   U�/V  pW�/V  0Yjustforfun_justforfun_ �/V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �|��O �u; /      Some_stuffs P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �n���O w�; /      Meeting /V  ���/V   ��/V  `�justforfun_justforfun_ �/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  ���?��O �^< /      Birthday    ��/V  `�/V  �#Some_stuffs_Some_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P�S��O :�I /      Appointment  U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  `ZA��O LiJ /      Birthday    P�/V  PQ�/V  0HThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  ���<��O G�V /      Birthday V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ���{��O �W /      Meeting     0s�/V  pt�/V  �uThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  0]�Ǯ�O N@W /      Appointment �Z�/V  �[�/V  �RSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   j���O ��Z /      Some_stuffs � �/V  0�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  0a����O >}f /      Workout /V  �	�/V  �/V  PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �V�P��O �uj /       Workout     P�/V  PQ�/V  0Hjustforfun_justforfun_ �/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V   *����O \�u /      Birthday    0]�/V  p^�/V  �_This_stuffs_This_stuffs_ /V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  h(7��O �5v /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �Z����O ��w /      Appointment P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  @Rx��O X�w /      Some_stuffs  <�/V  �F�/V  @?Some_stuffs_Some_stuffs_ /V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  ��.<��O Fd� /      Workout /V  ���/V  0��/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  @      h=�L��O 5�� /      Meeting /V  � �/V  0�/V  pThis_stuffs_This_stuffs_ /V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  �FA3�O �� /   	   Workout     P�/V  PQ�/V  0HSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  ����O �_� /       Appointment ���/V   ��/V  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V  ��*��O �-� /      Appointment ��/V  p�/V  pThis_stuffs_This_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  �<��O *̕ /      Meeting     ��/V   �/V  p+This_stuffs_This_stuffs_ /V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �C	>�O 㲖 /      Meeting     м�/V  ��/V  @�This_stuffs_This_stuffs_ /V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  h����O � /   	   Appointment  ��/V  @��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  �xaU�O �W� /       Meeting /V  P 
�/V  �
�/V  
This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  
�/V  �$
�/V  �%
�/V   
�/V  `
�/V  �
�/V  
�/V  P
�/V  �
�/V  P
�/V  �
�/V  �
�/V  
�/V  P
�/V  � 
�/V  "
�/V  :
�/V   '
�/V  `(
�/V  �)
�/V  �*
�/V   ,
�/V  �-
�/V   /
�/V  `0
�/V  �1
�/V  �8C��O �� /      Workout     ��/V  `�/V  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V   �&}/�O 8>� /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             @�}�1�O ��� /      Workout     ���/V   ��/V  `�This_stuffs_This_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  ���X3�O f�� /      Appointment ���/V   ��/V  `�This_stuffs_This_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  �(��L�O �� /      Workout     `��/V  ���/V  0�justforfun_justforfun_ �/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  XJ��N�O K�� /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��O�O �$� /      Meeting     �Z�/V  �[�/V  �RSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V  �.��Y� /      Birthday V  �9Կ&V   ;Կ&V  �<�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �GԿ&V  `IԿ&V  �PԿ&V   LԿ&V  @MԿ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  �.��Y@� /      Birthday V   RԿ&V  �SԿ&V   U�justforfun_justforfun_ Կ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  pԿ&V  �xԿ&V  �yԿ&V  p{Կ&V  �|Կ&V  ��Կ&V   �Կ&V  ��Կ&V  �.��Y� /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �.��Y� /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �.��Y@� /      Birthday    �	�/V  �/V  Pjustforfun_justforfun_ �/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  !m4�n�� /       Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               "m4�n�$� /      Some_stuffs ��/V  p�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  #m4�n�� /       Some_stuffs Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  �g��SW� /      Workout      ��/V  @��/V  ��Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  pI�*�3� /      Workout      ��/V  ���/V  ��justforfun_justforfun_ �/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �a����F^v /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �a����F]q /      Some_stuffs  ��/V  @��/V  ��Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  �a����F^v /      Birthday V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ��7�!S�. /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ��7�!S�2 /      Appointment ���/V  ���/V   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  ��7�!S�. /      Workout     Ј�/V  P��/V  ЏSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  �����u,	�"+ /      Meeting      <�/V  �F�/V  @?justforfun_justforfun_ �/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  �'/�)<	�+ /      Workout     @3	�/V  �4	�/V  �5	justforfun_justforfun_ 	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �t8n�Ah	�r- /      Some_stuffs ��/V  `�/V  �#Some_stuffs_Some_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  Y��&\��
9 /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             Z��&\��
K9 /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             [��&\��
9 /      Birthday V   <�/V  �F�/V  @?Some_stuffs_Some_stuffs_ /V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  !E�H]7�
q�; /      Some_stuffs `FԿ&V  �GԿ&V  `I�justforfun_justforfun_ Կ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  "E�H]7�
$�; /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     #E�H]7�
q�; /      Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               !���]�x�G /      Appointment  RԿ&V  �SԿ&V   U�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  pԿ&V  �xԿ&V  �yԿ&V  p{Կ&V  �|Կ&V  ��Կ&V   �Կ&V  ��Կ&V  "���]�D�G /      Appointment � �/V  0�/V  pSome_stuffs_Some_stuffs_ /V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  #���]�x�G /      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     A\�^*��H /   	   Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     A\�^* �H /      Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             A\�^*��H /   	   Meeting     P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �-ap,x�K /       Some_stuffs  �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �-ap,x<�K /       Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �-ap,x�K /       Some_stuffs ��/V  p�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  �8�&���W /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �8�&�� X /      Appointment ���/V  ���/V  �justforfun_justforfun_ �/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  �8�&���W /      Meeting     p��/V  ���/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  �w�5c���X /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �w�5c���X /   	   Some_stuffs  U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �w�5c���X /      Some_stuffs ���/V   ��/V  ��Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  Q�؃�J�X /      Workout     P�/V  PQ�/V  0HSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  R�؃���X /      Appointment  <�/V  �F�/V  @?Some_stuffs_Some_stuffs_ /V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  S�؃�5�X /      Appointment P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �瞴03�[ /      Some_stuffs ��/V  `�/V  �justforfun_justforfun_ �/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  �瞴037[ /      Appointment P�/V  PQ�/V  0HSome_stuffs_Some_stuffs_ /V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  �瞴03~[ /   	   Meeting     0��/V  ���/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V  AnC� �f /   	   Meeting     �ӿ&V  p�ӿ&V  p��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  P�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  BnC� �
f /      Birthday    ���/V  ���/V   �Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  CnC� �f /   	   Meeting     ���/V  `��/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  ���՞.x�f /   	   Some_stuffs  k	�/V  `l	�/V  �\	Some_stuffs_Some_stuffs_ /V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V   �	�/V  @�	�/V  )�.�>$^Mwh /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             *�.�>$^%|h /      Workout     ���/V  ���/V   �Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  +�.�>$^Mwh /      Meeting /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  i�ڰYj��h /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             j�ڰYj�h /      Birthday    Ј�/V  P��/V  ЏSome_stuffs_Some_stuffs_ /V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  k�ڰYj��h /      Meeting /V  �z�/V  ���/V  �~This_stuffs_This_stuffs_ /V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Qˊ���ow /      Some_stuffs ��/V  p�/V  pSome_stuffs_Some_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  ����`5�8�w /      Appointment P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V   ����dx� /      Appointment Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  _���ԓ /   	   Appointment  �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  _���Г /      Workout     ���/V  @��/V  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  _���ԓ /   	   Appointment ��/V  `�/V  �#This_stuffs_This_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  �,��UT4�� /      Some_stuffs PIӿ&V  �Jӿ&V  �M�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �,��UT~�� /      Appointment @��/V  ���/V  `�Some_stuffs_Some_stuffs_ /V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  `��/V  0��/V  p��/V  ���/V   ��/V  `��/V  �,��UT4�� /      Some_stuffs Ј�/V  P��/V  ЏThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  �ᒲ��d'� /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �ᒲ��d�(� /       Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               �ᒲ��d'� /      Birthday    P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  I����=lQo� /      Workout &V   �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  J����=lIu� /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             K����=lQo� /      Workout /V  ���/V  P��/V  �Some_stuffs_Some_stuffs_ /V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V  p���s /      Workout     ��/V  p�/V  pThis_stuffs_This_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  �j�*˘w�� /      Birthday V  ��/V  P��/V  ��This_stuffs_This_stuffs_ /V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  �j�*˘w7� /      Workout     ��/V  p�/V  pThis_stuffs_This_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  �j�*˘w�� /      Meeting     P|	�/V  �}	�/V  �m	Some_stuffs_Some_stuffs_ /V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  H�y�WN��� /      Meeting /V  �Q	�/V  �R	�/V  T	Some_stuffs_Some_stuffs_ /V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  ЕlŻ<��X� /      Birthday    �#�/V  P%�/V  �)Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  a��'�lٳ /      Some_stuffs p��/V  ���/V  ��This_stuffs_This_stuffs_ /V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �/V  P�/V  b��'��۳ /      Birthday    ��/V  p�/V  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  c��'��ڳ /      Some_stuffs Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  �Iǚ1K� /      Some_stuffs  �ҿ&V  p�ҿ&V  0��justforfun_justforfun_ ҿ&V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �Iǚ1��� /      Some_stuffs P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �Iǚ1K� /      Some_stuffs  U�/V  pW�/V  0Yjustforfun_justforfun_ �/V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  !�u�m.�}
 /      Appointment �z�/V  ���/V  �~This_stuffs_This_stuffs_ /V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  ��(~�m.k�
 /      Some_stuffs ���/V  ���/V  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V  0~��n.� /       Birthday    Ј�/V  P��/V  ЏThis_stuffs_This_stuffs_ /V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  �5U�n.k) /      Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ���J�n.�O /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             9�_��n.� /      Appointment �	�/V  P�	�/V  ��	This_stuffs_This_stuffs_ /V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  Ю	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ���(Ko.� /      Appointment �T
�/V  pV
�/V  �W
This_stuffs_This_stuffs_ /V  �]
�/V  0_
�/V  p`
�/V  �a
�/V  �z
�/V  �{
�/V  Pf
�/V  �g
�/V  i
�/V  Pj
�/V  �k
�/V  �l
�/V  n
�/V  Po
�/V  �p
�/V  Pr
�/V  �s
�/V  u
�/V  �v
�/V  �w
�/V  y
�/V  �
�/V  0}
�/V  p~
�/V  �
�/V  ��
�/V  0�
�/V  p�
�/V  ��
�/V  ��B�o.5� /   	   Some_stuffs ���/V  ���/V   �This_stuffs_This_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  ��C� p.�* /      Birthday V  PZ	�/V  �[	�/V  `L	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  F�p.4N /      Workout     p��/V  0��/V  ��Some_stuffs_Some_stuffs_ /V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  �n�ax.�� /      Meeting     � �/V  0�/V  pjustforfun_justforfun_ �/V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  �~�Ēx.f /      Workout /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  Qo���x.� /      Meeting /V  ��	�/V  0�	�/V  p�	justforfun_justforfun_ 	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  �
�/V  �
�/V  ��	�/V  �	�/V  P 
�/V  �
�/V  
�/V  P
�/V  �
�/V  
�/V  �
�/V  

�/V  �
�/V  
�/V  �$
�/V  �%
�/V   
�/V  `
�/V  �
�/V  
�/V  P
�/V  �
�/V  P
�/V  8����y.�� /      Workout     ��/V  p�/V  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  �-�Дz.K( /      Appointment  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ��aȂ.��* /      Appointment  U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  h�!��.M+ /      Birthday    �	�/V  0�	�/V  p�	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  0�	�/V  p�	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  p�	�/V  @�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  �^hz�.ڙ+ /       Some_stuffs � �/V  0�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  `�s߭�.��+ /      Birthday    P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �����.�[, /      Birthday    Ј�/V  P��/V  ЏThis_stuffs_This_stuffs_ /V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  �vb�1�.�, /      Birthday    ��/V  `�/V  �Some_stuffs_Some_stuffs_ /V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  Ph���.�B- /      Some_stuffs ���/V  ���/V   �Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  ����+�./�8 /      Appointment 0]�/V  p^�/V  �_justforfun_justforfun_ �/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  	�����.*�9 /      Workout     0]�/V  p^�/V  �_This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  C&L�.�: /       Birthday     ��/V  @��/V  ��This_stuffs_This_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  �U�tC�.�c: /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             a�7���.�u; /      Appointment `��/V  ��/V  `�This_stuffs_This_stuffs_ /V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  `��/V  0��/V  p��/V  ���/V   ��/V  `��/V  ���/V  0��/V  �)��.��; /      Appointment ���/V  Д�/V  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ()�Ub�.E< /       Workout /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  k����.�f< /      Some_stuffs  <�/V  �F�/V  @?This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  �����.��H /      Some_stuffs Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  P��Y-�.J_I /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �1mw�.��I /       Some_stuffs ��/V  p�/V  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  a�2\ݗ.poJ /      Appointment �
�/V  
�/V  P
justforfun_justforfun_ 
�/V  �
�/V  
�/V  P
�/V  � 
�/V  "
�/V  :
�/V   '
�/V  `(
�/V  �)
�/V  �*
�/V   ,
�/V  �-
�/V   /
�/V  `0
�/V  �1
�/V  `3
�/V  �4
�/V   6
�/V  �7
�/V  �N
�/V  P;
�/V  �<
�/V  >
�/V  �?
�/V  A
�/V  PB
�/V  �C
�/V  �D
�/V  F
�/V  �ogx�.�SK /       Workout     �$	�/V   &	�/V  `'	Some_stuffs_Some_stuffs_ /V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  9�U&�.��V /      Birthday    Ј�/V  P��/V  ЏThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  9w�>�.�W /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             q��H\�.-AW /      Some_stuffs ���/V   ��/V  @�Some_stuffs_Some_stuffs_ /V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V   �<ŧ�.d�W /      Appointment P$�/V  �%�/V   'This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  P����.�Y /   	   Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �I���.��Y /      Appointment �z�/V  ���/V  �~justforfun_justforfun_ �/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  ���1G�.>&Z /      Workout     �	�/V  �/V  PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  U ^�.�HZ /      Appointment �#�/V  P%�/V  �)This_stuffs_This_stuffs_ /V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  ���`��._�Z /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ��:Ţ.��Z /      Meeting     �R�/V  �S�/V  UThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  �	�=�./f /      Meeting     0s�/V  pt�/V  �uThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  �0�iq�.{}f /      Workout /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ���ť�.\�f /      Workout     ��	�/V  П	�/V  `�	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  Ю	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V   ����.�lg /      Workout /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  H���>�.ɳg /      Workout     ��/V  p�/V  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  ��1���.�h /       Some_stuffs `M�/V  �N�/V  �ZThis_stuffs_This_stuffs_ /V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  �`>�.�yj /      Appointment ��	�/V  0�	�/V  p�	Some_stuffs_Some_stuffs_ /V  ��	�/V  P�	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  0�	�/V  ��	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  �
�/V  �
�/V  ��	�/V  �	�/V  P 
�/V  �
�/V  
�/V  P
�/V  �
�/V  
�/V  �
�/V  

�/V  �
�/V  
�/V  �$
�/V  �K�ˣ�.��u /      Meeting     ��	�/V  Щ	�/V  �	justforfun_justforfun_ 	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  �Pش.�8v /       Birthday    p��/V  ��/V  0�This_stuffs_This_stuffs_ /V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  p�/V  p�/V  x���?�.o�v /       Workout     Ј�/V  P��/V  ЏThis_stuffs_This_stuffs_ /V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  (�p���.EEw /      Appointment @@	�/V  �A	�/V  �B	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  ��µ.0�w /   	   Appointment ���/V  0��/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  ��_7��.q�w /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             H$�m�.�x /      Workout /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  8q��t�.�x /      Birthday    ��/V  p�/V  pSome_stuffs_Some_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  1^{�:�.e� /      Appointment ���/V  ���/V   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  �+���.��� /       Meeting /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �Ŭ�>�.u� /   	   Workout /V  �	�/V  �/V  PSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  +i��.W� /       Birthday    PZ	�/V  �[	�/V  `L	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  (���.\_� /      Workout /V  �c
�/V  e
�/V  �O
This_stuffs_This_stuffs_ /V  �T
�/V  pV
�/V  �W
�/V  pY
�/V  �Z
�/V  0\
�/V  �]
�/V  0_
�/V  p`
�/V  �a
�/V  �z
�/V  �{
�/V  Pf
�/V  �g
�/V  i
�/V  Pj
�/V  �k
�/V  �l
�/V  n
�/V  Po
�/V  �p
�/V  Pr
�/V  �s
�/V  u
�/V  �v
�/V  �w
�/V  y
�/V  �
�/V  0}
�/V  ��
 ��.�� /      Workout     ���/V  @��/V  p�Some_stuffs_Some_stuffs_ /V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  X�n���.�m� /      Some_stuffs  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �x#V�.n1� /      Meeting     P�/V  PQ�/V  0HSome_stuffs_Some_stuffs_ /V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  Q��ܾ�.
ʕ /      Appointment @��/V  � 	�/V  �	This_stuffs_This_stuffs_ /V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  .I�W�.8�� /      Some_stuffs `��/V  ���/V  0�justforfun_justforfun_ �/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  �N����.� /      Birthday V  ��	�/V   �	�/V  @�	Some_stuffs_Some_stuffs_ /V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V   �	�/V  `�	�/V  ��	�/V  P�	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  0�	�/V  ��	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  �
�/V  �
�/V  ��	�/V  �	�/V  P 
�/V  �+B���.XR� /       Appointment ���/V   ��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  Q�Kt@�.�� /       Workout     P�/V  ��/V  This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �a�\�.p=� /      Birthday    ���/V  ���/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  ���`��.�>� /      Meeting     ���/V  Ъ�/V  P�justforfun_justforfun_ �/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V  ��,8��.��� /       Some_stuffs Ј�/V  P��/V  ЏSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  1W�@&�.�� /      Workout /V  �C
�/V  �D
�/V  F
Some_stuffs_Some_stuffs_ /V  K
�/V  �L
�/V  �c
�/V  e
�/V  �O
�/V  0Q
�/V  pR
�/V  �S
�/V  �T
�/V  pV
�/V  �W
�/V  pY
�/V  �Z
�/V  0\
�/V  �]
�/V  0_
�/V  p`
�/V  �a
�/V  �z
�/V  �{
�/V  Pf
�/V  �g
�/V  i
�/V  Pj
�/V  �k
�/V  �l
�/V  n
�/V  Po
�/V  �p
�/V  Xٝ���.Kx� /      Birthday    ��/V  `�/V  �#This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  ؈o"��.{�� /   	   Workout     p��/V  ���/V  ��Some_stuffs_Some_stuffs_ /V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �/V  P�/V  A9��"�.7�� /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               0��>�.�Ǵ /      Birthday    P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  Y�q���.1�� /      Some_stuffs ��/V  p�/V  pThis_stuffs_This_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  ���%�.�)� /      Appointment 0s�/V  pt�/V  �uThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  �B9�?y%Pz� /      Workout     P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V   ���#.$� /      Some_stuffs ��ӿ&V  P�ӿ&V  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  1z�ι�#.) /   	   Appointment ���/V  ���/V  �Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  2z�ι�#.n /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �$\n��#.�S /       Appointment @��/V  ���/V  ��Some_stuffs_Some_stuffs_ /V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @      �$\n��#.�O /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �4Z�l$.$� /      Birthday V  P�/V  ��/V  justforfun_justforfun_ �/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �4Z�l$.5� /   	   Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �ݷ	lx$.�& /      Birthday    `�/V  ��/V  �	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �ݷ	lx$.p' /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               ���$.]q /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��V�'.�� /      Birthday    ��	�/V  0�	�/V  p�	Some_stuffs_Some_stuffs_ /V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  �
�/V  �
�/V  ��	�/V  �	�/V  P 
�/V  �
�/V  
�/V  P
�/V  �
�/V  
�/V  �
�/V  

�/V  �
�/V  
�/V  �$
�/V  �%
�/V   
�/V  `
�/V  �
�/V  
�/V  P
�/V  �
�/V  P
�/V  ��V�'.'� /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ���)�(.2 /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     9�"G�J(.� /      Workout      ��/V  @��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  :�"G�J(.�� /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �^��[�+.q�* /       Meeting     P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �^��[�+.��* /      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     i69�+.� + /      Workout     ��/V  0��/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  j69�+.�+ /   	   Meeting /V  ��	�/V  ��	�/V   �	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  a��� (,.v�+ /      Workout      ��/V  @��/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  b��� (,.��+ /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��
F,.(^, /      Some_stuffs  U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ��
F,.�[, /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             Q$p!��,.rK- /      Birthday     ��/V  `��/V  мSome_stuffs_Some_stuffs_ /V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  R$p!��,.�G- /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             X3��a�/.K9 /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��:vo�/.�f: /      Appointment �	�/V  �/V  PSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  ��:vo�/.�c: /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                              Eo�EA0.$�; /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ))K}V0.�< /      Workout     P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  *)K}V0.�< /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                      һօi3.D�G /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             Ɍ���3.��H /      Workout     ���/V   ��/V  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  `��/V  0��/V  p��/V  ���/V  ʌ���3.��H /      Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                                ��.�3. �H /      Appointment ��ӿ&V  p�ӿ&V  0��This_stuffs_This_stuffs_ &V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  Q�/��3.YI /      Birthday V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  R�/��3.J_I /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �;�G4.�XK /   	   Meeting     ���/V  Ъ�/V  P�justforfun_justforfun_ �/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V  �;�G4.�TK /       Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �m� e4.<�K /       Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               !+@b�y7.Y�W /       Appointment @@	�/V  �A	�/V  �B	justforfun_justforfun_ 	�/V  �G	�/V  0I	�/V  PZ	�/V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  "+@b�y7.ɯW /       Workout &V  p[ӿ&V  �\ӿ&V  0`�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  �� ��7.� X /      Appointment  �ҿ&V  p�ҿ&V  0��justforfun_justforfun_ ҿ&V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �_T��7.�X /   	   Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     P@Q���7.J�X /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     Q�b�7. Y /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             R�b�7.�Y /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �1�U �7.`�Y /      Appointment ���/V  P��/V  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V  �1�U �7.��Y /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               �#���8.�'Z /      Appointment ��/V   �/V  �!This_stuffs_This_stuffs_ /V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  �#���8.>&Z /      Workout &V  �6Կ&V  `8Կ&V   >�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   BԿ&V  @CԿ&V  �JԿ&V  `FԿ&V  �GԿ&V  `IԿ&V  �PԿ&V   LԿ&V  @MԿ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @      ���$8.MZ /      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ���$8.cGZ /      Appointment  �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �ó;�98.��Z /       Birthday V  ��/V  P��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  �ó;�98._�Z /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ��bEX8.�[ /      Some_stuffs p[ӿ&V  �\ӿ&V  0`�justforfun_justforfun_ ӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  @~�Z�.;.�
f /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��C/8;.�1f /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ��C/8;.Q1f /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �&���`;. �f /      Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �&���`;.>�f /      Workout &V  p[ӿ&V  �\ӿ&V  0`�justforfun_justforfun_ ӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  !is�D�;.Hhg /       Meeting /V   <�/V  �F�/V  @?Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  "is�D�;.�lg /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             I�����;.��g /      Appointment ���/V  0��/V  p�justforfun_justforfun_ �/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  J�����;.ɳg /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     (L3
q�;.%|h /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��� o�;.��h /      Meeting /V  @��/V  ���/V  ��Some_stuffs_Some_stuffs_ /V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  ��� o�;.�h /       Some_stuffs ��ӿ&V  p�ӿ&V  0��This_stuffs_This_stuffs_ &V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  h#�.��;.�h /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             y<P��?.��v /      Appointment ���/V  0��/V  p�Some_stuffs_Some_stuffs_ /V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  z<P��?.o�v /       Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             )�AĢ?.,Kw /   	   Appointment  U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  *�AĢ?.�Hw /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             I��U�?.Bx /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     J��U�?.�x /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     9`hc��?.�x /      Workout     ���/V  @��/V  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  :`hc��?.�x /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �Ƥ֔lC.6� /      Birthday     ��/V  @��/V  ��justforfun_justforfun_ �/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  �Ƥ֔lC.u� /   	   Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �����D.m�� /   	   Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �����D.�� /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             M�G.�Г /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     Y�&�,G.�i� /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               Z�&�,G.�m� /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �
�B(H.:;� /      Birthday V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �
�B(H.p=� /      Birthday    ��ӿ&V  P�ӿ&V  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  ���kK.~�� /      Appointment PIӿ&V  �Jӿ&V  �M�Some_stuffs_Some_stuffs_ &V  �Vӿ&V  @Xӿ&V  p[ӿ&V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �=���<K.�(� /       Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               HA��PK.Iu� /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��D[�mK.�� /      Birthday V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  Y�ή��N.�|� /      Some_stuffs ��/V  `�/V  �justforfun_justforfun_ �/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  Z�ή��N.Kx� /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ���1�BO.ݵ� /       Appointment ���/V  P��/V  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V  ���1�BO.{�� /   	   Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             `?�3KO.lٳ /      Some_stuffs ��ӿ&V  P�ӿ&V  ���This_stuffs_This_stuffs_ &V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  1�%ձ�O.CŴ /      Some_stuffs ���/V   ��/V  `�Some_stuffs_Some_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  2�%ձ�O.�Ǵ /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �	q��O.��� /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     !�n��s�9�r� /      Meeting     ���/V  ���/V  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  "�n��s�9#q� /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     #�n��s�9dx� /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               $�n��s�9�r� /      Meeting &V   �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  Y��oi�?E�� /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               Z��oi�?�� /       Appointment ��/V  p�/V  pSome_stuffs_Some_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  [��oi�?E�� /      Workout     `M�/V  �N�/V  �Zjustforfun_justforfun_ �/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  \��oi�?)�� /   	   Some_stuffs `��/V  ���/V  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  ]��oi�?��� /      Meeting     �		�/V  �
	�/V  	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  =��M޲L�(� /      Some_stuffs ���/V   ��/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V  =��M޲L�(� /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     =��M޲L�"� /       Meeting &V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  =��M޲L�(� /      Some_stuffs  �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  =��M޲L�+� /      Some_stuffs ���/V  ���/V   �Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  =��M޲L�(� /      Meeting     P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V   =uɊܯR�+� /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             @�YSȥ /       Birthday V  �	�/V  P	�/V  �		This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �Eˣ`�YR� /      Meeting     ��/V  `�/V  �#Some_stuffs_Some_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  �Eˣ`�Y�� /      Some_stuffs ��ӿ&V  p�ӿ&V  0��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  �Eˣ`�YW� /      Workout &V  PIӿ&V  �Jӿ&V  �M�Some_stuffs_Some_stuffs_ &V  �Vӿ&V  @Xӿ&V  p[ӿ&V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �Eˣ`�YR� /      Meeting &V   �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  q�c�fa&a߽� /   	   Birthday V  ��
�/V  ��
�/V  0�
This_stuffs_This_stuffs_ /V  ��
�/V   �
�/V  `�
�/V  ��
�/V  ��
�/V   �
�/V  P�
�/V  ��
�/V  Е
�/V  P�
�/V  ��
�/V  Й
�/V  �
�/V  ��
�/V  �
�/V  ��
�/V  Р
�/V  �
�/V  p�
�/V  ��
�/V  �
�/V  0�
�/V  @�
�/V  ��
�/V  @�
�/V  ��
�/V   �
�/V  @�
�/V  ��
�/V  r�c�fa&a��� /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             s�c�fa&aN�� /       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     t�c�fa&a��� /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             q���}L"l� /      Appointment ���/V  0��/V  p�Some_stuffs_Some_stuffs_ /V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  r���}L"l� /      Meeting &V   �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  s���}L"l/� /   	   Some_stuffs p[ӿ&V  �\ӿ&V  0`�Some_stuffs_Some_stuffs_ &V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  t���}L"l� /      Meeting /V   ��/V  `��/V  мSome_stuffs_Some_stuffs_ /V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  A�oi��l9� /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             B�oi��l�� /   	   Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     C�oi��l� /   	   Appointment  �ҿ&V  p�ҿ&V  0��justforfun_justforfun_ ҿ&V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  D�oi��lȥ /       Birthday    PIӿ&V  �Jӿ&V  �M�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  E�oi��l9� /      Some_stuffs ��/V  p�/V  pThis_stuffs_This_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  F�oi��l�� /   	   Workout     ���/V  ���/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  G�oi��l� /   	   Appointment ��/V  p�/V  pjustforfun_justforfun_ �/V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  Iڗ3KR�vF� /      Birthday    P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  Jڗ3KR�v�� /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               Kڗ3KR�vK� /      Appointment ��ӿ&V  p�ӿ&V  0��This_stuffs_This_stuffs_ &V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  Lڗ3KR�v�� /      Birthday    ���/V  @��/V  p�justforfun_justforfun_ �/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  Y�5�]x� /      Birthday V  �ӿ&V  p�ӿ&V  p��justforfun_justforfun_ ӿ&V  �ӿ&V  `�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  �PMe�^�$+ /      Workout     �0	�/V   2	�/V  @3	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �PMe�^�%+ /   	   Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �PMe�^�a#+ /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �PMe�^�%+ /   	   Meeting /V   <�/V  �F�/V  @?Some_stuffs_Some_stuffs_ /V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  	1�	�����nw /   	   Some_stuffs ��/V  p�/V  pjustforfun_justforfun_ �/V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  
1�	����-mw /       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     1�	�����ow /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             1�	�����nw /   	   Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               �A��푵�,�w /      Workout /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �A��푵�C�w /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �A��푵���w /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �A��푵�C�w /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �7N����ͼ+ /      Meeting     ��	�/V  Ж	�/V  �	Some_stuffs_Some_stuffs_ /V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  Ю	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  �7N����"�+ /      Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �7N����"�+ /   	   Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �7N����"�+ /      Appointment  ��/V  @��/V  ��This_stuffs_This_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  �����̥�x� /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �����̥/}� /   	   Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �����̥�z� /       Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �����̥Pz� /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �����̥/}� /   	   Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �D��f��Wq- /      Meeting     p��/V  P��/V  ��This_stuffs_This_stuffs_ /V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  �D��f���r- /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               �D��f���r- /      Some_stuffs  �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �D��f��Wq- /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             XP�HU���� /       Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��pq��*X� /      Workout     0H�/V  pI�/V  �JSome_stuffs_Some_stuffs_ /V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  ��pq��GT� /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ��pq��W� /       Workout &V  `IԿ&V  �PԿ&V   L�justforfun_justforfun_ Կ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  pԿ&V  �xԿ&V  ��pq��GT� /      Birthday V  ��/V  `�/V  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  �.X��6��f /      Birthday     �	�/V  `�	�/V  ��	justforfun_justforfun_ 	�/V  p�	�/V  ��	�/V  0�	�/V  ��	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  �
�/V  �
�/V  ��	�/V  �	�/V  P 
�/V  �
�/V  
�/V  P
�/V  �
�/V  
�/V  �
�/V  

�/V  �
�/V  
�/V  �$
�/V  �%
�/V   
�/V  `
�/V  �
�/V  �.X��6f /       Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �.X��6�ȣf /      Appointment p[ӿ&V  �\ӿ&V  0`�justforfun_justforfun_ ӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  �.X��6f /       Appointment ���/V   ��/V  `�Some_stuffs_Some_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  