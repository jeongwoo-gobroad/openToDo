ܦ
 /   ��
 /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �< /   �< /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             8{ /   H{ /      Meeting                        This_stuffs_                                                                                                                                                                                                                                                         | /   � /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �lw /   -mw /       Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ,q /   ]q /      Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         \�; /   w�; /      Meeting                        justforfun                                                                                                                                                                                                                                                           }f /   >}f /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �c: /   �c: /      Workout                        This_stuffs_                                                                                                                                                                                                                                                         �|� /   /}� /   	   Workout                        This_stuffs_                                                                                                                                                                                                                                                         P� /   h� /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �G- /   �G- /      Meeting                        This_stuffs_                                                                                                                                                                                                                                                         � /   9� /      Some_stuffs                    This_stuffs_                                                                                                                                                                                                                                                         ��H /   ��H /      Some_stuffs                    justforfun                                                                                                                                                                                                                                                           l+� /   �+� /      Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         �p� /   #q� /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �= /   �= /      Meeting                        This_stuffs_                                                                                                                                                                                                                                                          9 /   K9 /      Workout                        This_stuffs_                                                                                                                                                                                                                                                         4�V /   G�V /      Birthday                       This_stuffs_                                                                                                                                                                                                                                                         �Ǵ /   �Ǵ /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             4� /   g� /       Birthday                       justforfun                                                                                                                                                                                                                                                           D�v /   o�v /       Workout                        This_stuffs_                                                                                                                                                                                                                                                         �y /   (�y /      Workout                        justforfun                                                                                                                                                                                                                                                           X' /   p' /      Birthday                       justforfun                                                                                                                                                                                                                                                           ;< /   A;< /      Birthday                       justforfun                                                                                                                                                                                                                                                           � /   '� /      Appointment                    Some_stuffs_                                                                                                                                                                                                                                                         -q /   ^v /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �|� /   �z� /       Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         �z� /   �z� /       Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ؓ� /   ٓ� /       Some_stuffs                    This_stuffs_                                                                                                                                                                                                                                                         lqZ /   uqZ /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             t� /   u� /   	   Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��� /   ��� /      Birthday                       Some_stuffs_                                                                                                                                                                                                                                                         <�f /   \�f /      Workout                        justforfun                                                                                                                                                                                                                                                           �X /   �X /   	   Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             P� /   }� /       Some_stuffs                    justforfun                                                                                                                                                                                                                                                           N� /   $N� /      Appointment                    justforfun                                                                                                                                                                                                                                                           �[, /   �[, /      Birthday                       This_stuffs_                                                                                                                                                                                                                                                         ��J /   ��J /   	   Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��
 /   ��
 /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �r+ /   s+ /      Workout �U   �e�U  p�e�U  0�eThis_stuffs_This_stuffs_ �U   f�U  �f�U  �f�U   f�U  f�U  �f�U  �f�U   f�U  @f�U  �f�U  f�U  �f�U  �f�U  Pf�U  �f�U   !f�U  �#f�U  �$f�U  �&f�U  p(f�U   ,f�U  �-f�U  0f�U  �2f�U  @5f�U  �6f�U  p9f�U  �:f�U  �=f�U  �;i /   �;i /      Workout                        Some_stuffs_                                                                                                                                                                                                                                                         ��� /   N�� /       Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �Г /   �Г /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             \D� /   fD� /      Meeting                        justforfun                                                                                                                                                                                                                                                            �+ /   "�+ /      Appointment                    This_stuffs_                                                                                                                                                                                                                                                         �Ǵ /   CŴ /      Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         @T� /   GT� /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �*� /   �*� /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             _I /   J_I /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �TK /   �TK /       Appointment                    This_stuffs_                                                                                                                                                                                                                                                         du; /   �u; /      Some_stuffs                    justforfun                                                                                                                                                                                                                                                           h� /   �� /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             `H+ /   wH+ /   	   Some_stuffs                    justforfun                                                                                                                                                                                                                                                           4� /   5� /   	   Some_stuffs                    This_stuffs_                                                                                                                                                                                                                                                         ��Z /   ��Z /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             8�w /   X�w /      Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         �(� /   �(� /       Some_stuffs                    justforfun                                                                                                                                                                                                                                                           xlg /   �lg /      Workout                        Some_stuffs_                                                                                                                                                                                                                                                         �|� /   Pz� /      Workout                        This_stuffs_                                                                                                                                                                                                                                                         �lw /   �ow /      Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         8؆ /   V؆ /      Appointment                    justforfun                                                                                                                                                                                                                                                           �1 /   2 /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             4�� /   5�� /      Meeting                        This_stuffs_                                                                                                                                                                                                                                                         !9 /   9 /      Birthday                       Some_stuffs_                                                                                                                                                                                                                                                         4� /   :� /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �x /   �x /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��� /   ��� /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �lw /   �nw /   	   Some_stuffs                    justforfun                                                                                                                                                                                                                                                           �X /   �X /      Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         H�� /   {�� /   	   Workout                        Some_stuffs_                                                                                                                                                                                                                                                         |?� /   ~?� /      Meeting                        justforfun                                                                                                                                                                                                                                                           `MX /   `MX /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             u� /   Iu� /      Meeting                        Some_stuffs_                                                                                                                                                                                                                                                         �: /   �: /      Birthday                       justforfun                                                                                                                                                                                                                                                           m+� /   �(� /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �Y /   �Y /      Workout                        This_stuffs_                                                                                                                                                                                                                                                         <~
 /   d~
 /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �� /   �� /      Workout                        justforfun                                                                                                                                                                                                                                                           5� /   $� /      Birthday                       justforfun                                                                                                                                                                                                                                                           <@W /   N@W /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �x /   Bx /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��� /   ��� /      Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         �, /   9�, /       Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �-� /   �-� /      Appointment                    This_stuffs_                                                                                                                                                                                                                                                         �1 /   . /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             � /   � /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �c: /   �f: /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��* /   ��* /      Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         d� /   Fd� /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             xO /   �O /      Workout                        This_stuffs_                                                                                                                                                                                                                                                         �r- /   �r- /      Appointment                    justforfun                                                                                                                                                                                                                                                           �m� /   �m� /      Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         \�+ /   ��+ /      Birthday                       This_stuffs_                                                                                                                                                                                                                                                         ��g /   ɳg /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �p� /   dx� /      Appointment                    justforfun                                                                                                                                                                                                                                                           �{h /   %|h /      Workout                        Some_stuffs_                                                                                                                                                                                                                                                         �G /   D�G /      Appointment                    Some_stuffs_                                                                                                                                                                                                                                                         �$+ /   %+ /   	   Meeting                        Some_stuffs_                                                                                                                                                                                                                                                         ��, /   ��, /       Meeting                        This_stuffs_                                                                                                                                                                                                                                                          �; /   $�; /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                              �K /   <�K /       Birthday                       justforfun                                                                                                                                                                                                                                                           �+ /   "�+ /   	   Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             d� /   �� /      Birthday                       justforfun                                                                                                                                                                                                                                                           0x� /   Kx� /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             u� /   6� /      Birthday                       justforfun                                                                                                                                                                                                                                                           � /   �� /   	   Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �˕ /   *̕ /      Meeting                        This_stuffs_                                                                                                                                                                                                                                                         ��� /   ʷ� /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��g /   ��g /      Appointment                    justforfun                                                                                                                                                                                                                                                           Ԕ� /   Ք� /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             D�Z /   _�Z /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             TPu /   �Pu /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �(� /   '� /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ࡗ /   �� /       Appointment                    Some_stuffs_                                                                                                                                                                                                                                                         �h /   �h /      Birthday                       Some_stuffs_                                                                                                                                                                                                                                                         �
f /   �
f /      Birthday                       Some_stuffs_                                                                                                                                                                                                                                                         P�K /   _�K /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ylg /   Hhg /       Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �$+ /   a#+ /      Meeting                        Some_stuffs_                                                                                                                                                                                                                                                         �m� /   �i� /      Workout                        justforfun                                                                                                                                                                                                                                                           �[ /   �[ /   	   Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �{h /   Mwh /      Meeting                        Some_stuffs_                                                                                                                                                                                                                                                         �?8 /   �?8 /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ̌W /   όW /       Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �� /   �� /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��f /   ��f /       Appointment                    Some_stuffs_                                                                                                                                                                                                                                                         8}x /   :}x /      Meeting                        This_stuffs_                                                                                                                                                                                                                                                         �� /   P�� /   	   Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��Y /   ��Y /      Appointment                    justforfun                                                                                                                                                                                                                                                           ��Y /   `�Y /      Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             @�w /   C�w /      Birthday                       justforfun                                                                                                                                                                                                                                                           ��� /   K� /      Some_stuffs  �e�U  p�e�U  0�ejustforfun   ��e�U  �e�U   f�U  �f�U  �f�U   f�U  f�U  �f�U  �f�U   f�U  @f�U  �f�U  f�U  �f�U  �f�U  Pf�U  �f�U   !f�U  �#f�U  �$f�U  �&f�U  p(f�U   ,f�U  �-f�U  0f�U  �2f�U  @5f�U  �6f�U  p9f�U  �:f�U  �=f�U  ha� /   ha� /      Meeting �U  PIf�U  �Jf�U  �MfThis_stuffs_This_stuffs_ �U  �Vf�U  @Xf�U  p[f�U  �\f�U  0`f�U  �af�U   ef�U  �ff�U  �if�U  `kf�U  �nf�U  �of�U  Psf�U  �tf�U  `xf�U  �yf�U  @}f�U  �~f�U  p�f�U  ��f�U  0�f�U  ��f�U  ��f�U   �f�U  ��f�U  `�f�U  �f�U  ��f�U  ��f�U  � /   6� /      Workout �U  ��f�U  P�f�U  ��fjustforfun   ��f�U   �f�U  ��f�U  @�f�U  ��f�U  p�f�U  0�f�U  p�f�U  @�f�U  ��f�U  `�f�U  ��f�U  ��f�U  �f�U  ��f�U  P�f�U  `g�U  �g�U  �g�U  @	g�U  pg�U  �g�U  0g�U  pg�U  �g�U  �g�U   "g�U  `#g�U  �(g�U  P*g�U  �/g�U  ]�+ /   v�+ /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �p� /   �r� /      Meeting �U   �e�U  p�e�U  0�eSome_stuffs_Some_stuffs_ �U   f�U  �f�U  �f�U   f�U  f�U  �f�U  �f�U   f�U  @f�U  �f�U  f�U  �f�U  �f�U  Pf�U  �f�U   !f�U  �#f�U  �$f�U  �&f�U  p(f�U   ,f�U  �-f�U  0f�U  �2f�U  @5f�U  �6f�U  p9f�U  �:f�U  �=f�U  1x� /   �|� /      Some_stuffs PIf�U  �Jf�U  �Mfjustforfun    Rf�U  �Sf�U  �Vf�U  @Xf�U  p[f�U  �\f�U  0`f�U  �af�U   ef�U  �ff�U  �if�U  `kf�U  �nf�U  �of�U  Psf�U  �tf�U  `xf�U  �yf�U  @}f�U  �~f�U  p�f�U  ��f�U  0�f�U  ��f�U  ��f�U   �f�U  ��f�U  `�f�U  �f�U  ��f�U  ��f�U  �&X /   �&X /      Birthday U  �f�U  p�f�U  p�fSome_stuffs_  �f�U  ��f�U  �f�U  `�f�U  ��f�U  P�f�U  ��f�U  P�f�U  ��f�U   �f�U  ��f�U  @�f�U  ��f�U  p�f�U  0�f�U  p�f�U  @�f�U  ��f�U  `�f�U  ��f�U  ��f�U  �f�U  ��f�U  P�f�U  `g�U  �g�U  �g�U  @	g�U  pg�U  �g�U  0g�U  L /   n /      Meeting                        This_stuffs_                                                                                                                                                                                                                                                         � X /   � X /      Appointment  �e�U  p�e�U  0�ejustforfun   ��e�U  �e�U   f�U  �f�U  �f�U   f�U  f�U  �f�U  �f�U   f�U  @f�U  �f�U  f�U  �f�U  �f�U  Pf�U  �f�U   !f�U  �#f�U  �$f�U  �&f�U  p(f�U   ,f�U  �-f�U  0f�U  �2f�U  @5f�U  �6f�U  p9f�U  �:f�U  �=f�U  ,�f /   >�f /      Workout �U  p[f�U  �\f�U  0`fjustforfun    ef�U  �ff�U  �if�U  `kf�U  �nf�U  �of�U  Psf�U  �tf�U  `xf�U  �yf�U  @}f�U  �~f�U  p�f�U  ��f�U  0�f�U  ��f�U  ��f�U   �f�U  ��f�U  `�f�U  �f�U  ��f�U  ��f�U  �f�U  �f�U  `�f�U  @�f�U  ��f�U  �f�U  p�f�U  p�f�U  ��� /   ��� /   	   Appointment ��f�U  p�f�U  0�fSome_stuffs_Some_stuffs_ �U  `�f�U  ��f�U  ��f�U  �f�U  ��f�U  P�f�U  `g�U  �g�U  �g�U  @	g�U  pg�U  �g�U  0g�U  pg�U  �g�U  �g�U   "g�U  `#g�U  �(g�U  P*g�U  �/g�U  P1g�U  �6g�U  `8g�U   >g�U  @?g�U  �9g�U   ;g�U  �<g�U  \�; /   ��; /      Workout                        Some_stuffs_                                                                                                                                                                                                                                                         !�K /   �K /       Some_stuffs  �e�U  p�e�U  0�eThis_stuffs_This_stuffs_ �U   f�U  �f�U  �f�U   f�U  f�U  �f�U  �f�U   f�U  @f�U  �f�U  f�U  �f�U  �f�U  Pf�U  �f�U   !f�U  �#f�U  �$f�U  �&f�U  p(f�U   ,f�U  �-f�U  0f�U  �2f�U  @5f�U  �6f�U  p9f�U  �:f�U  �=f�U  �� /   � /   	   Appointment PIf�U  �Jf�U  �MfThis_stuffs_This_stuffs_ �U  �Vf�U  @Xf�U  p[f�U  �\f�U  0`f�U  �af�U   ef�U  �ff�U  �if�U  `kf�U  �nf�U  �of�U  Psf�U  �tf�U  `xf�U  �yf�U  @}f�U  �~f�U  p�f�U  ��f�U  0�f�U  ��f�U  ��f�U   �f�U  ��f�U  `�f�U  �f�U  ��f�U  ��f�U  p' /   �' /      Meeting �U  ��f�U  P�f�U  ��fThis_stuffs_ ��f�U   �f�U  ��f�U  @�f�U  ��f�U  p�f�U  0�f�U  p�f�U  @�f�U  ��f�U  `�f�U  ��f�U  ��f�U  �f�U  ��f�U  P�f�U  `g�U  �g�U  �g�U  @	g�U  pg�U  �g�U  0g�U  pg�U  �g�U  �g�U   "g�U  `#g�U  �(g�U  P*g�U  �/g�U  D�) /   J�) /      Meeting                        justforfun                                                                                                                                                                                                                                                           �uj /   �uj /       Workout �U   �e�U  p�e�U  0�ejustforfun   ��e�U  �e�U   f�U  �f�U  �f�U   f�U  f�U  �f�U  �f�U   f�U  @f�U  �f�U  f�U  �f�U  �f�U  Pf�U  �f�U   !f�U  �#f�U  �$f�U  �&f�U  p(f�U   ,f�U  �-f�U  0f�U  �2f�U  @5f�U  �6f�U  p9f�U  �:f�U  �=f�U  ��u /   ��u /      Some_stuffs p[f�U  �\f�U  0`fThis_stuffs_This_stuffs_ �U  �if�U  `kf�U  �nf�U  �of�U  Psf�U  �tf�U  `xf�U  �yf�U  @}f�U  �~f�U  p�f�U  ��f�U  0�f�U  ��f�U  ��f�U   �f�U  ��f�U  `�f�U  �f�U  ��f�U  ��f�U  �f�U  �f�U  `�f�U  @�f�U  ��f�U  �f�U  p�f�U  p�f�U  