                                                                �g����  ��/      Workout     �x��fU  py��fU  0}�cillum dolore eu fugiat nulla pariatur ��fU  ���fU  Ћ��fU  �����  ��/       Birthday    �z��fU  �{��fU  `|�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �����  ��/       Birthday    `���fU   ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �����  ��/       Birthday     Q��fU  �Q��fU  U�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �����  ��/       Birthday    ���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��S���  e/      Birthday nt 0
��fU  �
��fU  0�cillum dolore eu fugiat nulla pariatur roident ��fU   ��fU  ������  �3/       Workout     ��fU  ���fU  P�cillum dolore eu fugiat nulla pariatur ��fU  ��fU  ���fU  ������  �3/       Workout  ion i��fU  �i��fU   j�cillum dolore eu fugiat nulla pariatur im id est laborum. U  ������  �3/       Workout  ion k��fU  �k��fU  Pl�cillum dolore eu fugiat nulla pariatur im id est laborum. U  ������  �3/       Workout  ion u��fU  �u��fU  v�cillum dolore eu fugiat nulla pariatur im id est laborum. U  $�����  84/      Meeting     �&��fU  p'��fU  �)�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  @�|���  h_/       consectetur ����fU  ����fU  P��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   A�|���  h_/       consectetur @���fU  ����fU  @��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �c����  ��/       bonorum fU  �s��fU  pt��fU  0u�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �c����  ��/       bonorum tion T��fU   U��fU  �U�Lorem ipsum dolor sit amet, consectetur adipiscing elit .    �c����  ��/       bonorum tion ��fU   ��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit .    �c����  ��/       bonorum tion W��fU  �W��fU  pX�Lorem ipsum dolor sit amet, consectetur adipiscing elit .    �w����  ��/      exercitation ���fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  �37���  ��/      Appointment  ���fU  ���fU  `��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �o����  -�/       consectetur P��fU   ��fU  P�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �o����  -�/       consectetur ^��fU  �^��fU  _�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �����  �/      consectetur `j��fU  �j��fU  �v�Duis aute irure dolor in rehendert in volupate velit esse U  pGe���  /       Appointment @���fU   ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  qGe���  /       Appointment ���fU  `���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  rGe���  /       Appointment ���fU  ��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  sGe���  /       Appointment ���fU  0��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  ����  5J/       Meeting     ����fU  @���fU  ���cillum dolore eu fugiat nulla pariatur ��fU   ���fU  ����fU  	����  5J/       Meeting     �1��fU  �2��fU  `3�cillum dolore eu fugiat nulla pariatur ��fU  �7��fU  `8��fU  ����  $p/      malorum     �d��fU  `e��fU   f�Duis aute irure dolor in rehendert in volupate velit esse U  �I����  H�/      malorum     p��fU  0��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Խi���  ��/      bonorum fU  B��fU  pL��fU  �C�Duis aute irure dolor in rehendert in volupate velit esse U  yw���  J�/       bonorum     ���fU  @ ��fU  � �ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  yw���  J�/       bonorum     @f��fU   g��fU  �j�ullamco laboris nisi ut aliquip ex ea commodo consequat e U  ����  _0/       Birthday     6��fU  �6��fU  �7�Excepteur sint occaecat cupidatat non proident ��fU  �<��fU  ����  _0/       Birthday                       Excepteur sint occaecat cupidatat non proident               ����  _0/       Birthday    @���fU  ����fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  ����  _0/       Birthday    `���fU   ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU   ���fU  \����  �0/      Meeting     D��fU  �D��fU  �G�cillum dolore eu fugiat nulla pariatur ��fU  U��fU  �U��fU  ������  �/      Workout     ���fU  `��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �9k���  è/       Birthday    0���fU  ����fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �9k���  è/       Birthday nt  q��fU  �q��fU  `r�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �	���  /�/      exercitation ��fU  P��fU  �Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  x$����  ��/       bonorum     @f��fU   g��fU  �j�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   z$����  ��/       bonorum tion ���fU  `���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   |$����  ��/       bonorum tion ���fU  `���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   $����  ��/       bonorum tion *��fU   +��fU  �+�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ~q����  �/       Workout     `���fU   ���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �q����  �/       Workout tur  ���fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat iq   �Ч���  ��/       consectetur P��fU  ���fU  � �sunt in culpa qui offici desunt molit aim id est laborum. U  �Ч���  ��/       consectetur P���fU  ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  �Ч���  ��/       consectetur p���fU  ����fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  �Ч���  ��/       consectetur  ��fU  ���fU  `�sunt in culpa qui offici desunt molit aim id est laborum. U  ��+���  �/      Workout                        cillum dolore eu fugiat nulla pariatur                       ��,���  �/       Birthday    @���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ��,���  �/       Birthday    �z��fU  {��fU  �{�Duis aute irure dolor in rehendert in volupate velit esse U  ��5���  $/       Birthday                       Excepteur sint occaecat cupidatat non proident               ��5���  $/       Birthday    ���fU  `��fU   �Excepteur sint occaecat cupidatat non proident ��fU  �$��fU  ��5���  $/       Birthday    p���fU  0���fU  ��Excepteur sint occaecat cupidatat non proident ��fU  p���fU  ��5���  $/       Birthday    pm��fU   n��fU  �n�Excepteur sint occaecat cupidatat non proident ��fU  Pr��fU  �%����  pF/       Appointment                    sunt in culpa qui offici desunt molit aim id est laborum.    �%����  pF/       Appointment P5��fU  �5��fU  P6�sunt in culpa qui offici desunt molit aim id est laborum. U  �%����  pF/       Appointment ?��fU  �?��fU  �@�sunt in culpa qui offici desunt molit aim id est laborum. U  �%����  pF/       Appointment �M��fU  N��fU  �N�sunt in culpa qui offici desunt molit aim id est laborum. U  ��j���  4m/      bonorum     �&��fU  p'��fU  �)�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  H�����  ]�/       exercitation                   Lorem ipsum dolor sit amet, consectetur adipiscing elit      I�����  ]�/       exercitation ���fU  `���fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  J�����  ]�/       exercitation ���fU  `���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  K�����  ]�/       exercitation ���fU  ����fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  Qp$���  R�/       Appointment ����fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  Sp$���  R�/       Appointment `���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  Up$���  R�/       Appointment p���fU  ����fU  p��Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  Wp$���  R�/       Appointment @���fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  H55���  ��/       malorum fU  P��fU  ��fU  `�sunt in culpa qui offici desunt molit aim id est laborum. U  J55���  ��/       malorum     P���fU  ���fU  p��sunt in culpa qui offici desunt molit aim id est laborum. U  L55���  ��/       malorum     `3��fU   4��fU  �4�sunt in culpa qui offici desunt molit aim id est laborum. U  N55���  ��/       malorum     g��fU  �g��fU  Ph�sunt in culpa qui offici desunt molit aim id est laborum. U  )"����  i/       exercitation ��fU  0��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  *"����  i/       exercitation +��fU  �+��fU  0,�Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   d�����  @/      Birthday    �&��fU  p'��fU  �)�sunt in culpa qui offici desunt molit aim id est laborum. U  <����  W�#/      Appointment �A��fU  PB��fU  �B�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �#��  �#/       bonorum     ���fU  p���fU  0��sunt in culpa qui offici desunt molit aim id est laborum. U  �#��  �#/       bonorum tion p��fU  pq��fU  @��sunt in culpa qui offici desunt molit aim id est laborum. U  ̓-��  ��#/      Appointment                    sed do eiusmo tempo incidunt ut labore et dolor magna aliq   \�;��  �'$/      consectetur ����fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��@��  #)$/       exercitation ���fU  ���fU  ���Excepteur sint occaecat cupidatat non proident onsequat �fU  ��@��  #)$/       exercitation ���fU  `���fU  ��Excepteur sint occaecat cupidatat non proident onsequat �fU  qPR��  �-$/       Birthday    @f��fU   g��fU  �j�cillum dolore eu fugiat nulla pariatur ��fU  �x��fU  py��fU  tPR��  �-$/       Birthday    ���fU  ����fU  ��cillum dolore eu fugiat nulla pariatur ��fU  0���fU  ����fU  �eU��  p.$/       malorum fU  �{��fU   |��fU  �|�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �eU��  p.$/       malorum     ���fU  p���fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �b���  $/      bonorum     `3��fU   4��fU  �4�sunt in culpa qui offici desunt molit aim id est laborum. U  !� ��  �$/       bonorum     ����fU  p���fU  0��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  #� ��  �$/       bonorum     ����fU  `���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �,!��  $�$/       Meeting     ���fU  `��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  �,!��  $�$/       Meeting  nt ��fU  ���fU  P�Duis aute irure dolor in rehendert in volupate velit esse U  ����  9�$/       exercitation ���fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  ����  9�$/       exercitation ���fU   ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ����  9�$/       exercitation ���fU  P���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  ����  9�$/       exercitation ��fU  `��fU   �Duis aute irure dolor in rehendert in volupate velit esse U  �bJ ��  :�$/      consectetur ���fU  p��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  ��� ��  :%/      Birthday                       cillum dolore eu fugiat nulla pariatur                       q6h!��  f9%/       malorum                        Lorem ipsum dolor sit amet, consectetur adipiscing elit      s6h!��  f9%/       malorum fU  ����fU  @���fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  u6h!��  f9%/       malorum     0J��fU  �J��fU  0K�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  w6h!��  f9%/       malorum      T��fU  �T��fU  0U�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  P�x!��  �=%/       malorum                        ullamco laboris nisi ut aliquip ex ea commodo consequat      R�x!��  �=%/       malorum     ����fU   ���fU  P��ullamco laboris nisi ut aliquip ex ea commodo consequat e U  T�x!��  �=%/       malorum     ����fU  ����fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat e U  V�x!��  �=%/       malorum     p���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat e U  d
�"��  @�%/      Meeting     @���fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  �=#��  ��%/      Meeting fU  p^��fU  0_��fU  �_�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �8�#��  y�%/       exercitation |��fU  `}��fU  �}�sunt in culpa qui offici desunt molit aim id est laborum. U  �8�#��  y�%/       exercitation ��fU  ���fU  `�sunt in culpa qui offici desunt molit aim id est laborum. U  `<
%��  |'&/       malorum     ��fU  ���fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  a<
%��  |'&/       malorum     ���fU  0��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  ���%��  Q&/      Workout                        sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �?&��  �v&/      exercitation ��fU  �!��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  <�`'��  ��&/      Workout     l��fU  �l��fU  m�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  $	�'��  ��&/      Birthday    @���fU   ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  �9�(��  q'/      Workout fU  P,��fU  -��fU  �-�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   XG�(��  �'/       malorum                        ullamco laboris nisi ut aliquip ex ea commodo consequat      ZG�(��  �'/       malorum tur ����fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  [G�(��  �'/       malorum tur ����fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  \G�(��  �'/       malorum tur  ���fU  ����fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��1)��  �7'/      malorum fU  P���fU  ����fU  P��cillum dolore eu fugiat nulla pariatur ��fU  ���fU  н��fU  P�a*��  ��'/       exercitation ���fU  `���fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  Q�a*��  ��'/       exercitation ��fU  ���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  R�a*��  ��'/       exercitation ��fU  ���fU  P�Duis aute irure dolor in rehendert in volupate velit esse U  U�a*��  ��'/       exercitation ��fU  ���fU  P�Duis aute irure dolor in rehendert in volupate velit esse U  4�o*��  �'/       bonorum     ����fU  ����fU  0��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  6�o*��  �'/       bonorum ent  ��fU  ���fU  0�ullamco laboris nisi ut aliquip ex ea commodo consequat e U  O�r*��  �'/      malorum     ����fU  @���fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  ���*��  )�'/      Appointment  =��fU  �=��fU  `@�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  @^�*��  h�'/       Appointment                    sed do eiusmo tempo incidunt ut labore et dolor magna aliq   B^�*��  h�'/       Appointment `���fU  ����fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   C^�*��  h�'/       Appointment ����fU  P���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   D^�*��  h�'/       Appointment ���fU  P��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   4R�+��  B�'/      Appointment Ш��fU  ����fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��+W��  ��2/      Workout     ����fU  `���fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  p�W��  �3/       Appointment  R��fU  �R��fU   S�cillum dolore eu fugiat nulla pariatur ��fU   W��fU  �W��fU  p�W��  �3/       Appointment �L��fU  M��fU  �M�cillum dolore eu fugiat nulla pariatur ��fU  �P��fU  PQ��fU  ظ�W��  w!3/       consectetur p(��fU  0)��fU  0*�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ٸ�W��  w!3/       consectetur 0��fU  ���fU  0�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ڸ�W��  w!3/       consectetur �I��fU  @J��fU  �J�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ݸ�W��  w!3/       consectetur  0��fU  �0��fU  01�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  B�W��  �$3/      Workout     p���fU  0���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU  P���fU  ��CX��  �D3/      Birthday    P���fU  ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �KX��  �F3/       Birthday    P���fU  ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �KX��  �F3/       Birthday    `���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �KX��  �F3/       Birthday    �v��fU  `w��fU  �w�Duis aute irure dolor in rehendert in volupate velit esse U  �KX��  �F3/       Birthday    ���fU  ����fU  P��Duis aute irure dolor in rehendert in volupate velit esse U  ���Y��  G�3/      Meeting     `3��fU   4��fU  �4�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �q
Z��  �3/      Workout      ���fU  ����fU  @��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��Z��  ��3/       consectetur 0���fU  ����fU  p��sunt in culpa qui offici desunt molit aim id est laborum. U  ��Z��  ��3/       consectetur ���fU  �	��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  ��Z��  ��3/       consectetur  ���fU  ����fU   ��sunt in culpa qui offici desunt molit aim id est laborum. U  ��Z��  ��3/       consectetur  ���fU  ����fU  `��sunt in culpa qui offici desunt molit aim id est laborum. U  0!�Z��  ��3/      malorum     0s��fU  �s��fU  �x�sunt in culpa qui offici desunt molit aim id est laborum. U  ��Z��  J�3/       Workout fU  �x��fU  py��fU  0}�Excepteur sint occaecat cupidatat non proident velit esse U  ��Z��  J�3/       Workout fU  `���fU   ���fU  ��Excepteur sint occaecat cupidatat non proident velit esse U  ��Z��  J�3/       Workout     ����fU  ����fU   ��Excepteur sint occaecat cupidatat non proident velit esse U  ��Z��  J�3/       Workout     ����fU  ����fU  `��Excepteur sint occaecat cupidatat non proident velit esse U  �l�Z��  v�3/       exercitation ��fU  0��fU  ��cillum dolore eu fugiat nulla pariatur ��fU  � ��fU  `!��fU  �l�Z��  v�3/       exercitation ���fU  ����fU   x�cillum dolore eu fugiat nulla pariatur ��fU  `|��fU  �|��fU  ��k\��  �T4/      consectetur D��fU  �D��fU  �G�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �¾]��  ��4/       Meeting     D��fU  �D��fU  �G�Excepteur sint occaecat cupidatat non proident ��fU  �U��fU  �¾]��  ��4/       Meeting     Ш��fU  ����fU  ��Excepteur sint occaecat cupidatat non proident velit esse U  �¾]��  ��4/       Meeting     ��fU  ���fU  P�Excepteur sint occaecat cupidatat non proident velit esse U  �¾]��  ��4/       Meeting      0��fU  �0��fU  P1�Excepteur sint occaecat cupidatat non proident velit esse U  ��4^��  ��4/       consectetur @f��fU   g��fU  �j�Excepteur sint occaecat cupidatat non proident ��fU  py��fU  ��4^��  ��4/       consectetur 0
��fU  �
��fU  0�Excepteur sint occaecat cupidatat non proident ��fU   ��fU  ��4^��  ��4/       consectetur  W��fU  �W��fU  `X�Excepteur sint occaecat cupidatat non proident ��fU  P]��fU  ��4^��  ��4/       consectetur  ���fU  ����fU  ���Excepteur sint occaecat cupidatat non proident ��fU   ���fU  '�B^��  x�4/      Birthday U  ����fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ���^��  ��4/      exercitation                   Lorem ipsum dolor sit amet, consectetur adipiscing elit      	��^��  ��4/       consectetur `���fU  ���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ���fU  ����fU  
��^��  ��4/       consectetur �&��fU  �'��fU  p(�cillum dolore eu fugiat nulla pariatur  adipiscing elit iq   $|�_��  �5/      Appointment �L��fU  �M��fU  pN�Duis aute irure dolor in rehendert in volupate velit esse U  �*`��  �A5/      bonorum     ����fU  `���fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  �``��  yE5/       Appointment B��fU  pL��fU  �C�cillum dolore eu fugiat nulla pariatur ��fU   H��fU  �H��fU  �``��  yE5/       Appointment @f��fU   g��fU  �j�cillum dolore eu fugiat nulla pariatur ��fU  �x��fU  py��fU  �``��  yE5/       Appointment ����fU  @���fU  ���cillum dolore eu fugiat nulla pariatur ��fU   ���fU  ����fU  �``��  yE5/       Appointment ����fU  `���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU  ����fU  <)�`��  wg5/      consectetur                    Excepteur sint occaecat cupidatat non proident               ĽBa��  �5/      malorum                        cillum dolore eu fugiat nulla pariatur                       ���a��  Q�5/      Appointment ����fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��gb��  �5/      malorum fU  �+��fU  p,��fU  �,�sunt in culpa qui offici desunt molit aim id est laborum. U  �lc��  S	6/      Meeting     �6��fU  `7��fU  �7�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   (�c��  �06/      Birthday    ���fU  ����fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  e\.d��  �Q6/      Workout     @f��fU   g��fU  �j�Excepteur sint occaecat cupidatat non proident ��fU  py��fU  ��;d��  �T6/       Appointment ����fU  ����fU  p��Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  ��;d��  �T6/       Appointment p��fU  ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  ��;d��  �T6/       Appointment ���fU  �	��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  ��;d��  �T6/       Appointment ����fU  ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  0��d��  �z6/       Birthday                       Duis aute irure dolor in rehendert in volupate velit esse    2��d��  �z6/       Birthday U  ����fU  p���fU  0��Duis aute irure dolor in rehendert in volupate velit esse U  3��d��  �z6/       Birthday    P���fU  О��fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  5��d��  �z6/       Birthday    ����fU  0���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ���d��  $|6/       Workout     ���fU  ���fU  �sunt in culpa qui offici desunt molit aim id est laborum. U  ���d��  $|6/       Workout     pj��fU  �j��fU  pk�sunt in culpa qui offici desunt molit aim id est laborum. U  %/�d��  �|6/      Birthday    P��fU  ��fU  `�Duis aute irure dolor in rehendert in volupate velit esse U  9^e��  J�6/       Birthday     g��fU  �g��fU   h�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   9^e��  J�6/       Birthday    ���fU  ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   P>	f��  �6/       Meeting ent ����fU  ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat e U  Q>	f��  �6/       Meeting ent �T��fU  `U��fU  �U�ullamco laboris nisi ut aliquip ex ea commodo consequat e U  ��f��  9�6/       Appointment @���fU  ����fU  @��cillum dolore eu fugiat nulla pariatur ��fU  @���fU  ����fU  ��f��  9�6/       Appointment ���fU  @��fU  ��cillum dolore eu fugiat nulla pariatur ��fU  �"��fU  p#��fU  |�Ag��  7/      bonorum     ����fU  0���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��i��  �7/       Workout                        sunt in culpa qui offici desunt molit aim id est laborum.    ��i��  �7/       Workout tion m��fU  `n��fU  �n�sunt in culpa qui offici desunt molit aim id est laborum.    ��i��  �7/       Workout tion ���fU  ����fU   ��sunt in culpa qui offici desunt molit aim id est laborum.    ��i��  �7/       Workout tion ���fU  ����fU  p��sunt in culpa qui offici desunt molit aim id est laborum.    vA���  �^B/       exercitation                   sed do eiusmo tempo incidunt ut labore et dolor magna aliq   	vA���  �^B/       exercitation 1��fU  �1��fU  �2�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   
vA���  �^B/       exercitation ���fU  P���fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   vA���  �^B/       exercitation /��fU  �0��fU  �9�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �I���  �`B/      exercitation H��fU  `I��fU  PJ�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �+ܓ��  0�B/      Birthday U  <��fU  �<��fU  �=�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �w���  /�B/       Appointment ���fU  Ћ��fU  Џ�sunt in culpa qui offici desunt molit aim id est laborum. U  �w���  /�B/       Appointment @���fU  ����fU  @��sunt in culpa qui offici desunt molit aim id est laborum. U  �w���  /�B/       Appointment p���fU  0���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  �w���  /�B/       Appointment ����fU  ����fU   ��sunt in culpa qui offici desunt molit aim id est laborum. U  �����  C C/       Meeting     p���fU  0���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  p���fU  0���fU  �����  C C/       Meeting     ����fU  ����fU   ��cillum dolore eu fugiat nulla pariatur olupate velit esse U  �����  C C/       Meeting     ����fU  @���fU  ���cillum dolore eu fugiat nulla pariatur olupate velit esse U  �����  C C/       Meeting     p���fU  ���fU  ���cillum dolore eu fugiat nulla pariatur olupate velit esse U  6Q;���  �!C/       consectetur �4��fU   5��fU  �5�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  :Q;���  �!C/       consectetur �3��fU  4��fU  �4�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �<���  
"C/       Meeting     �9��fU  P:��fU  �1�sunt in culpa qui offici desunt molit aim id est laborum. U  �<���  
"C/       Meeting     �y��fU   z��fU  �z�sunt in culpa qui offici desunt molit aim id est laborum. U  �<���  
"C/       Meeting     0���fU  ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  �<���  
"C/       Meeting      F��fU  �F��fU   G�sunt in culpa qui offici desunt molit aim id est laborum. U  � X���  �(C/       Birthday    � ��fU  0!��fU  �!�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  � X���  �(C/       Birthday ur �j��fU  `k��fU  l�ullamco laboris nisi ut aliquip ex ea commodo consequat . U  �]���  l*C/       Meeting     p���fU  0���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �]���  l*C/       Meeting     ���fU  ���fU  p�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �]���  l*C/       Meeting fU  0���fU  ����fU  0��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �]���  l*C/       Meeting     ���fU  p��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ����  pLC/      Appointment D��fU  �D��fU  �G�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �o���  hpC/      malorum     p[��fU  0\��fU  �\�Excepteur sint occaecat cupidatat non proident ��fU  `b��fU  �����  �D/       Workout fU  ����fU  `���fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �����  �D/       Workout ent ����fU  `���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �����  �D/       Workout ent �\��fU  P]��fU  ^�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �����  �D/       Workout ent Pq��fU  �q��fU  Pr�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   u����  *D/      malorum     ���fU  Ћ��fU  Џ�Excepteur sint occaecat cupidatat non proident ��fU  0���fU  ����  �D/       malorum     ����fU  @���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ����  �D/       malorum     �z��fU  �{��fU  p|�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �w���  D7D/      bonorum     `���fU   ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ��}���  �8D/       malorum      ��fU  �!��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��}���  �8D/       malorum     ����fU  ���fU  Ч�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��}���  �8D/       malorum fU  ����fU  @���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��}���  �8D/       malorum      ���fU  ����fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   1�����  ��D/       exercitation ���fU  ����fU  @��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   2�����  ��D/       exercitation ���fU  @���fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   3�����  ��D/       exercitation ��fU  0��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   5�����  ��D/       exercitation ���fU   ���fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   <S����  ��D/      Meeting                        sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �=����  A�D/       malorum     ����fU  p���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �=����  A�D/       malorum     �w��fU  �x��fU  �y�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �K���  ܮD/      exercitation x��fU  py��fU  0}�ullamco laboris nisi ut aliquip ex ea commodo consequat e U  $�ܜ��  8�D/      exercitation W��fU  �W��fU  0X�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �Ip���  ��D/       bonorum     p���fU  ����fU  p��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �Ip���  ��D/       bonorum     0T��fU  �T��fU  pU�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   eZy���  @�D/      bonorum fU  `���fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   XȀ���  '�D/       bonorum fU  ����fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ZȀ���  '�D/       bonorum     `���fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat . U  [Ȁ���  '�D/       bonorum     ����fU  ���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat . U  ]Ȁ���  '�D/       bonorum     0	��fU  �	��fU  0
�ullamco laboris nisi ut aliquip ex ea commodo consequat . U  `���  �#E/       Workout     ���fU  P��fU  �Duis aute irure dolor in rehendert in volupate velit esse U  a���  �#E/       Workout     �8��fU  P9��fU  �9�Duis aute irure dolor in rehendert in volupate velit esse U  b���  �#E/       Workout     =��fU  �=��fU  `>�Duis aute irure dolor in rehendert in volupate velit esse U  c���  �#E/       Workout     ����fU  P���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  򳜞��  �FE/       bonorum fU  P��fU  ��fU  ��Excepteur sint occaecat cupidatat non proident ��fU  P��fU  ������  �FE/       bonorum     �+��fU  PM��fU  �,�Excepteur sint occaecat cupidatat non proident velit esse U  ������  �FE/       bonorum     ���fU  0��fU  ��Excepteur sint occaecat cupidatat non proident velit esse U  ������  �FE/       bonorum     � ��fU  �)��fU  p"�Excepteur sint occaecat cupidatat non proident velit esse U  ������  �GE/      Meeting                        sunt in culpa qui offici desunt molit aim id est laborum.    �ӥ���  ,IE/       Workout     0G��fU  �G��fU  0H�Duis aute irure dolor in rehendert in volupate velit esse U  �ӥ���  ,IE/       Workout     �H��fU   I��fU  �I�Duis aute irure dolor in rehendert in volupate velit esse U  �ǩ���  /JE/       Workout     �+��fU  p,��fU  �,�sunt in culpa qui offici desunt molit aim id est laborum. U  �ǩ���  /JE/       Workout     ��fU  ���fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  �ǩ���  /JE/       Workout     ���fU   ��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  �ǩ���  /JE/       Workout     �T��fU   U��fU  �U�sunt in culpa qui offici desunt molit aim id est laborum. U  �SI���  sE/      exercitation ���fU  @���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��K���  �sE/       exercitation z��fU  �{��fU  `|�sunt in culpa qui offici desunt molit aim id est laborum. U  ��K���  �sE/       exercitation ���fU  `���fU  ��sunt in culpa qui offici desunt molit aim id est laborum.    ��K���  �sE/       exercitation ���fU   ��fU  ���sunt in culpa qui offici desunt molit aim id est laborum.    ��K���  �sE/       exercitation ���fU   ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum.    �#O���  �tE/       malorum fU  p%��fU  0&��fU  �&�Duis aute irure dolor in rehendert in volupate velit esse U  �#O���  �tE/       malorum tur 0*��fU  �*��fU  �+�Duis aute irure dolor in rehendert in volupate velit esse U  �#O���  �tE/       malorum tur ���fU  P��fU  �Duis aute irure dolor in rehendert in volupate velit esse U  �#O���  �tE/       malorum tur �$��fU  `%��fU  0&�Duis aute irure dolor in rehendert in volupate velit esse U  0�؟��  ��E/       malorum     pU��fU  �`��fU  0W�cillum dolore eu fugiat nulla pariatur ��fU  p[��fU  0\��fU  1�؟��  ��E/       malorum fU  �$��fU  p%��fU  �%�cillum dolore eu fugiat nulla pariatur ��fU  P)��fU   *��fU  2�؟��  ��E/       malorum     �v��fU  `w��fU   l�cillum dolore eu fugiat nulla pariatur ��fU  `p��fU   q��fU  3�؟��  ��E/       malorum     PJ��fU  �J��fU  PK�cillum dolore eu fugiat nulla pariatur ��fU  �N��fU  PO��fU  �~���  D�E/      malorum     ����fU  ����fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ����  ��E/      exercitation ��fU  ��fU  `�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �#0���  01F/       exercitation ���fU  ����fU  @��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �#0���  01F/       exercitation A��fU  @B��fU  �B�Excepteur sint occaecat cupidatat non proident ��fU  pF��fU  o����  �UF/       bonorum      G��fU  �G��fU  �H�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  o����  �UF/       bonorum     �C��fU  `D��fU  �D�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  "�ˢ��  YF/       bonorum      ���fU  ����fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU  ����fU  $�ˢ��  YF/       bonorum tion ���fU  ����fU  `��cillum dolore eu fugiat nulla pariatur et dolor magna aliq   =�֢��  �[F/      exercitation ���fU  0���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  0�z���  ޅF/       exercitation z��fU  �{��fU  `|�cillum dolore eu fugiat nulla pariatur ��fU  `���fU  ����fU  1�z���  ޅF/       exercitation &��fU  p'��fU  �)�cillum dolore eu fugiat nulla pariatur ��fU   5��fU  �5��fU  2�z���  ޅF/       exercitation ���fU  ���fU  п�cillum dolore eu fugiat nulla pariatur ��fU  ����fU  P���fU  3�z���  ޅF/       exercitation ���fU  ����fU  `��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  `���fU  �>����  ��F/       Meeting     Ќ��fU  P���fU  Ѝ�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �>����  ��F/       Meeting     ����fU  ����fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   46���  ¨F/      malorum      l��fU  �l��fU  �m�cillum dolore eu fugiat nulla pariatur ��fU  �q��fU  �r��fU  �+K���  �{Q/      Workout     ����fU  `���fU   ��sunt in culpa qui offici desunt molit aim id est laborum. U  \ku���  �Q/      Birthday U   H��fU  �H��fU  �I�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   D����  ��Q/       Meeting     `p��fU   q��fU  �q�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  F����  ��Q/       Meeting     0S��fU  �S��fU  �T�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  )	����  ��Q/       Appointment ����fU   ���fU  P��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  *	����  ��Q/       Appointment P��fU  ���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  +	����  ��Q/       Appointment p���fU  0���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  -	����  ��Q/       Appointment ���fU  0��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  (�*���  i�Q/       Birthday    0G��fU  �G��fU  0H�cillum dolore eu fugiat nulla pariatur olupate velit esse    )�*���  i�Q/       Birthday    @���fU   ���fU  ���cillum dolore eu fugiat nulla pariatur olupate velit esse    ������  DR/       Appointment                    Lorem ipsum dolor sit amet, consectetur adipiscing elit      ������  DR/       Appointment ����fU  P���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ������  DR/       Appointment 0��fU  ���fU  0�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ������  DR/       Appointment ����fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  %����  xR/      Meeting     �&��fU  p'��fU  �)�Excepteur sint occaecat cupidatat non proident ��fU  �5��fU  ������  lR/       Workout     ����fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  ������  lR/       Workout     ���fU  ��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  ������  lR/       Workout      	��fU  ��fU  P
�Duis aute irure dolor in rehendert in volupate velit esse U  ������  lR/       Workout     p���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �x���  Q�R/      Workout     �X��fU  pY��fU  0Z�Duis aute irure dolor in rehendert in volupate velit esse U  ����  ��R/      consectetur                    sunt in culpa qui offici desunt molit aim id est laborum.    de����   �R/      Meeting     @���fU   ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ��<���  ;S/      Workout     p%��fU  0&��fU  �&�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  H�����  )S/       Workout fU  ����fU  ����fU  @��Excepteur sint occaecat cupidatat non proident ��fU  `���fU  I�����  )S/       Workout      H��fU  �H��fU  �I�Excepteur sint occaecat cupidatat non proident ��fU  �M��fU  J�����  )S/       Workout     Pc��fU  �c��fU  �d�Excepteur sint occaecat cupidatat non proident ��fU  �h��fU  K�����  )S/       Workout     �#��fU  `$��fU  �$�Excepteur sint occaecat cupidatat non proident ��fU  �(��fU  ��u���  [QS/      Appointment `?��fU  @��fU  �@�Excepteur sint occaecat cupidatat non proident ��fU  pD��fU  2}���  @SS/       Meeting ent ���fU  �	��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  2}���  @SS/       Meeting ent ����fU  ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  $,���  �vS/       consectetur 0U��fU  �U��fU  0V�sunt in culpa qui offici desunt molit aim id est laborum. U  &,���  �vS/       consectetur  ���fU  ����fU  ��sunt in culpa qui offici desunt molit aim id est laborum.    !���  xS/       Appointment                    Excepteur sint occaecat cupidatat non proident               "���  xS/       Appointment  ���fU  P���fU  ���Excepteur sint occaecat cupidatat non proident velit esse U  #���  xS/       Appointment  i��fU  �i��fU  `j�Excepteur sint occaecat cupidatat non proident velit esse U  %���  xS/       Appointment  ���fU  p���fU  0��Excepteur sint occaecat cupidatat non proident velit esse U  tQ%���  J~S/      Appointment                    Excepteur sint occaecat cupidatat non proident               ԡ���  *�S/       malorum fU  ����fU   ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  `���fU  ԡ���  *�S/       malorum     0���fU  Н��fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �����  ��S/       Meeting     P���fU  ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �����  ��S/       Meeting     � ��fU  P!��fU  �!�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �����  ��S/       Meeting     P��fU  ���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �����  ��S/       Meeting     :��fU  �:��fU  ;�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  6C����  �S/      Meeting                        sed do eiusmo tempo incidunt ut labore et dolor magna aliq   hk����  ��S/       Birthday    �n��fU  �o��fU  `p�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  kk����  ��S/       Birthday     ���fU  ����fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat . U  mk����  ��S/       Birthday    p���fU  ����fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat . U  pk����  ��S/       Birthday    ����fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat . U  6;���  n�S/      Workout     �&��fU  p'��fU  �)�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��T���  ��S/       consectetur                    Excepteur sint occaecat cupidatat non proident onsequat      ��T���  ��S/       consectetur =��fU  �=��fU  `>�Excepteur sint occaecat cupidatat non proident onsequat �fU  ��T���  ��S/       consectetur �6��fU  `7��fU  �7�Excepteur sint occaecat cupidatat non proident onsequat �fU  ��T���  ��S/       consectetur �7��fU  `8��fU   9�Excepteur sint occaecat cupidatat non proident onsequat �fU  ������  ��S/       exercitation D��fU  �D��fU  �G�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ������  ��S/       exercitation ��fU   ��fU  P�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ������  ��S/       exercitation ���fU  ����fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ������  ��S/       exercitation ���fU  0���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �����  (?T/      bonorum      
��fU  �
��fU  0�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �eL���  p�T/       Meeting      H��fU  �H��fU  �I�Excepteur sint occaecat cupidatat non proident ��fU  �M��fU  �eL���  p�T/       Meeting     0/��fU  �/��fU  ��Excepteur sint occaecat cupidatat non proident t laborum. U  �eL���  p�T/       Meeting fU  �	��fU  0
��fU  �
�Excepteur sint occaecat cupidatat non proident t laborum. U  �eL���  p�T/       Meeting      R��fU  �R��fU   S�Excepteur sint occaecat cupidatat non proident t laborum. U  ��l���  E�T/      consectetur U��fU  �U��fU  Y�cillum dolore eu fugiat nulla pariatur ��fU  @f��fU   g��fU  �\w���  ��T/       Workout  ion ���fU  p���fU  ��cillum dolore eu fugiat nulla pariatur  adipiscing elit �fU  �\w���  ��T/       Workout  ion F��fU  `G��fU  �G�cillum dolore eu fugiat nulla pariatur  adipiscing elit �fU  ������  C#U/       Appointment P1��fU  �1��fU  �2�Duis aute irure dolor in rehendert in volupate velit esse U  ������  C#U/       Appointment 0I��fU  �I��fU  0J�Duis aute irure dolor in rehendert in volupate velit esse U  ������  C#U/       Appointment �A��fU  PB��fU  �B�Duis aute irure dolor in rehendert in volupate velit esse U  ������  C#U/       Appointment p.��fU  0/��fU  �/�Duis aute irure dolor in rehendert in volupate velit esse U  ������  �'U/      Meeting     ����fU  @���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  �-���  %KU/      Workout      ���fU  ����fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �3���  �LU/       consectetur ���fU  `��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  �3���  �LU/       consectetur 0���fU  ����fU  0��Duis aute irure dolor in rehendert in volupate velit esse    �c���  �U/       exercitation s��fU  �s��fU  t�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �c���  �U/       exercitation ^��fU   _��fU  �_�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �]{���  ��U/      Birthday    U��fU  �U��fU  Y�sunt in culpa qui offici desunt molit aim id est laborum. U  ������  0�U/       consectetur �j��fU  �k��fU  l�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ������  0�U/       consectetur �]��fU  0^��fU  �^�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �v<���  �V/      Workout     ����fU  ����fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   D��	��  l�`/      Appointment @��fU   ��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  �,��  �a/      Appointment ���fU  P��fU  �Excepteur sint occaecat cupidatat non proident velit esse U  ����  :5a/       exercitation N��fU  PO��fU  �O�Excepteur sint occaecat cupidatat non proident ��fU  �S��fU  ����  :5a/       exercitation ���fU  ����fU  `��Excepteur sint occaecat cupidatat non proident velit esse U  7Y���  �6a/       Workout      
��fU  �
��fU  0�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ;Y���  �6a/       Workout     ��fU  ���fU  P�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �����  �7a/       Workout     ����fU  `���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �����  �7a/       Workout fU   ���fU  ����fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat e U  �����  �7a/       Workout     �^��fU  _��fU  �_�ullamco laboris nisi ut aliquip ex ea commodo consequat e U  �����  �7a/       Workout     l��fU  �l��fU  `m�ullamco laboris nisi ut aliquip ex ea commodo consequat e U  ����  �9a/       Appointment  6��fU  �6��fU  �7�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ����  �9a/       Appointment �4��fU  `5��fU   6�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ����  �9a/       Appointment  ��fU  ���fU   �Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ����  �9a/       Appointment �2��fU  3��fU  �3�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  9R��  �\a/       Workout      ���fU  ����fU  P��Excepteur sint occaecat cupidatat non proident ��fU  н��fU  :R��  �\a/       Workout fU  ����fU   ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  ,�_��  -`a/      exercitation ���fU  ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ����  �a/      malorum      ���fU  ����fU   ��sunt in culpa qui offici desunt molit aim id est laborum. U  m���  �a/      bonorum tur p���fU  ���fU   ��sunt in culpa qui offici desunt molit aim id est laborum.    ��!��  Y�a/       Appointment  ���fU  ����fU  `��sunt in culpa qui offici desunt molit aim id est laborum. U  ��!��  Y�a/       Appointment �,��fU  �-��fU  p.�sunt in culpa qui offici desunt molit aim id est laborum. U  ��!��  Y�a/       Appointment P1��fU  �1��fU  P2�sunt in culpa qui offici desunt molit aim id est laborum. U  ��!��  Y�a/       Appointment `r��fU   s��fU  �s�sunt in culpa qui offici desunt molit aim id est laborum. U  |z���  ��a/      Appointment p[��fU  0\��fU  �\�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ,	T��  �!b/      Appointment  H��fU  �H��fU  �I�cillum dolore eu fugiat nulla pariatur ��fU  �L��fU  �M��fU  y!Y��  #b/       Meeting fU  �^��fU   _��fU  �_�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   z!Y��  #b/       Meeting     ����fU  p���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   `���  \�b/       exercitation ��fU  ���fU  p�Excepteur sint occaecat cupidatat non proident onsequat �fU  b���  \�b/       exercitation P��fU  `Q��fU   R�Excepteur sint occaecat cupidatat non proident onsequat iq   d���  \�b/       exercitation ���fU  `���fU   ��Excepteur sint occaecat cupidatat non proident onsequat iq   g���  \�b/       exercitation ��fU  P ��fU  �"�Excepteur sint occaecat cupidatat non proident onsequat iq   Y����  '�b/       consectetur  ��fU  ���fU  ��cillum dolore eu fugiat nulla pariatur ��fU  ���fU  ���fU  [����  '�b/       consectetur                    cillum dolore eu fugiat nulla pariatur ommodo consequat      ]����  '�b/       consectetur  l��fU  �l��fU  `m�cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  `����  '�b/       consectetur  ���fU  `���fU   ��cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  rp���  վb/      consectetur ���fU  P��fU  �Excepteur sint occaecat cupidatat non proident ��fU   	��fU  !�<��  t�b/       malorum     ����fU  ����fU  `��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   #�<��  t�b/       malorum tur p(��fU  0)��fU  0*�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   %�<��  t�b/       malorum tur ���fU  @��fU   �sed do eiusmo tempo incidunt ut labore et dolor magna aliq   '�<��  t�b/       malorum tur P1��fU  �1��fU  �2�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��G��  M�b/       malorum     ����fU  ����fU   ��cillum dolore eu fugiat nulla pariatur ��fU  @���fU   ���fU  ��G��  M�b/       malorum     �&��fU  p'��fU  �)�cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  ��G��  M�b/       malorum     ����fU  P���fU  ���cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  ��G��  M�b/       malorum     ���fU  p���fU  ��cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  
'���  5c/       Meeting tur                    ullamco laboris nisi ut aliquip ex ea commodo consequat .    '���  5c/       Meeting tur ����fU  ����fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat . U  '���  5c/       Meeting tur ����fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat . U  '���  5c/       Meeting tur @���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat . U  ty���  Jc/      consectetur @���fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �����  �
c/       Appointment ���fU  Ћ��fU  Џ�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �����  �
c/       Appointment `���fU  ���fU  `��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �����  �
c/       Appointment �"��fU  p#��fU  �#�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �����  �
c/       Appointment �$��fU   %��fU  �%�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��r��  �/c/       malorum                        Duis aute irure dolor in rehendert in volupate velit esse    ��r��  �/c/       malorum     ����fU  P���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  ��r��  �/c/       malorum     n��fU  �n��fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ��r��  �/c/       malorum     `S��fU  0T��fU  �T�Duis aute irure dolor in rehendert in volupate velit esse U  �nt��  =0c/      Appointment P���fU  ���fU  У�sunt in culpa qui offici desunt molit aim id est laborum. U  d�B��  ��c/      bonorum     P��fU  ��fU  `�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �����  �c/       Meeting      H��fU  �H��fU  �I�Excepteur sint occaecat cupidatat non proident ��fU  �M��fU  �����  �c/       Meeting     P���fU  ����fU  ���Excepteur sint occaecat cupidatat non proident onsequat �fU  �����  �c/       Meeting  U  ����fU  ����fU  @��Excepteur sint occaecat cupidatat non proident onsequat �fU  �����  �c/       Meeting     p���fU   ���fU  ���Excepteur sint occaecat cupidatat non proident onsequat �fU   ����  ��c/       Meeting                        Excepteur sint occaecat cupidatat non proident               #����  ��c/       Meeting     �P��fU  `Q��fU   R�Excepteur sint occaecat cupidatat non proident velit esse U  &����  ��c/       Meeting fU  ����fU  ���fU  ���Excepteur sint occaecat cupidatat non proident velit esse U  )����  ��c/       Meeting     0Q��fU  �Q��fU  �R�Excepteur sint occaecat cupidatat non proident velit esse U  �����  ��c/       malorum                        ullamco laboris nisi ut aliquip ex ea commodo consequat      �����  ��c/       malorum fU  �4��fU  `5��fU  �5�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �����  ��c/       malorum     �'��fU  �(��fU  )�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ����  ��c/       malorum     �,��fU  �-��fU  p.�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �d��  ��c/      exercitation ���fU  ���fU  У�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �.��  �d/      Appointment ����fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  �z���  >Ed/      malorum fU  ����fU  ����fU  @��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  `���fU  ����  nFd/       Workout     P���fU  О��fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ����  nFd/       Workout     `q��fU  �q��fU  `r�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��5��  �gd/       Appointment ����fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  ��5��  �gd/       Appointment �O��fU  pP��fU  0Q�Duis aute irure dolor in rehendert in volupate velit esse U  ��5��  �gd/       Appointment ����fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  ��5��  �gd/       Appointment 0J��fU  �J��fU  0K�Duis aute irure dolor in rehendert in volupate velit esse U  �����  ��d/      Appointment ����fU  @���fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  �+���  ,�d/       consectetur `���fU   ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  �+���  ,�d/       consectetur ����fU  `���fU   ��sunt in culpa qui offici desunt molit aim id est laborum. U  �+���  ,�d/       consectetur  ���fU  ����fU   ��sunt in culpa qui offici desunt molit aim id est laborum. U  �+���  ,�d/       consectetur ����fU  `���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  �nw��  9�d/       Workout     `|��fU  �|��fU  �}�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �nw��  9�d/       Workout     P]��fU  �]��fU   y�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �_���  �e/       Workout fU   6��fU  �6��fU  �7�Excepteur sint occaecat cupidatat non proident ��fU  �<��fU  �_���  �e/       Workout     �-��fU  �.��fU  �C�Excepteur sint occaecat cupidatat non proident ing elit �fU  �_���  �e/       Workout      i��fU  �i��fU  `j�Excepteur sint occaecat cupidatat non proident ing elit �fU  �_���  �e/       Workout                        Excepteur sint occaecat cupidatat non proident ing elit      ����  te/      bonorum fU  �f��fU  `g��fU  �g�Excepteur sint occaecat cupidatat non proident onsequat �fU  U�wE��  ��o/      malorum fU  ����fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq    ��E��   p/       exercitation ��fU  p��fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��E��   p/       exercitation ���fU  ����fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  @5#F��  �)p/       Appointment                    Lorem ipsum dolor sit amet, consectetur adipiscing elit      B5#F��  �)p/       Appointment ���fU  `��fU   �Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  C5#F��  �)p/       Appointment  c��fU  �c��fU   d�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  D5#F��  �)p/       Appointment ����fU  P���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  m2F��  �-p/      Meeting     0���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  h��F��  QPp/       consectetur                    sed do eiusmo tempo incidunt ut labore et dolor magna aliq   j��F��  QPp/       consectetur P���fU  ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   k��F��  QPp/       consectetur �C��fU  @D��fU  00�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   l��F��  QPp/       consectetur 0J��fU  �J��fU  0K�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ~�F��  �Pp/      exercitation ���fU  ����fU  @��Excepteur sint occaecat cupidatat non proident ��fU  `���fU  � ]G��  %zp/      Meeting     @���fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �R�G��  >�p/      malorum                        cillum dolore eu fugiat nulla pariatur                       ��G��  ˠp/       bonorum     p���fU  0���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��G��  ˠp/       bonorum      ���fU  ����fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��G��  ˠp/       bonorum fU  @x��fU  �x��fU  �y�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��G��  ˠp/       bonorum     p���fU  ����fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��{H��  ��p/      bonorum fU   ���fU  ����fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  aI��  ��p/       Meeting tur `���fU   ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   cI��  ��p/       Meeting tur 0P��fU  �P��fU  0Q�Lorem ipsum dolor sit amet, consectetur adipiscing elit iq    �&I��  T�p/       Birthday    � ��fU  �)��fU  p"�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  "�&I��  T�p/       Birthday    ���fU  p��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  `'�I��  \q/       malorum                        sunt in culpa qui offici desunt molit aim id est laborum.    a'�I��  \q/       malorum  ur 0v��fU  �v��fU  pw�sunt in culpa qui offici desunt molit aim id est laborum. U  b'�I��  \q/       malorum  ur  ���fU  ����fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  c'�I��  \q/       malorum  ur 0���fU  ����fU  0��sunt in culpa qui offici desunt molit aim id est laborum. U  !�SJ��  T<q/       consectetur �9��fU  P:��fU  �1�Duis aute irure dolor in rehendert in volupate velit esse U  "�SJ��  T<q/       consectetur ����fU  @���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  #�SJ��  T<q/       consectetur ����fU  @���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  $�SJ��  T<q/       consectetur ����fU  ����fU  `��Duis aute irure dolor in rehendert in volupate velit esse U  ��XJ��  �=q/      consectetur p^��fU  0_��fU  �_�Duis aute irure dolor in rehendert in volupate velit esse U  x��J��  {aq/       Birthday U  ���fU  P��fU  �Excepteur sint occaecat cupidatat non proident ��fU  ���fU  y��J��  {aq/       Birthday    �q��fU  �r��fU  `s�Excepteur sint occaecat cupidatat non proident ing elit iq   z��J��  {aq/       Birthday    �&��fU  p'��fU  �)�Excepteur sint occaecat cupidatat non proident ing elit iq   {��J��  {aq/       Birthday    pj��fU  �j��fU  pk�Excepteur sint occaecat cupidatat non proident ing elit iq   ��K��  j�q/       Birthday     6��fU  �6��fU  �7�Duis aute irure dolor in rehendert in volupate velit esse U  ��K��  j�q/       Birthday    0Z��fU  �Z��fU  p[�Duis aute irure dolor in rehendert in volupate velit esse U  ��K��  j�q/       Birthday    V��fU  �V��fU  �L�Duis aute irure dolor in rehendert in volupate velit esse U  ��K��  j�q/       Birthday    �e��fU  Pf��fU  g�Duis aute irure dolor in rehendert in volupate velit esse U  �x�K��  ��q/       consectetur                    Lorem ipsum dolor sit amet, consectetur adipiscing elit      �x�K��  ��q/       consectetur ���fU  �	��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �x�K��  ��q/       consectetur ���fU  P��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �x�K��  ��q/       consectetur  ��fU  ���fU   �Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  `YL��  ��q/       consectetur P��fU  ��fU  `�cillum dolore eu fugiat nulla pariatur ��fU  �&��fU  p'��fU  cYL��  ��q/       consectetur ����fU  ����fU   ��cillum dolore eu fugiat nulla pariatur ��fU  @���fU   ���fU  eYL��  ��q/       consectetur ����fU  ���fU  ���cillum dolore eu fugiat nulla pariatur ��fU   ���fU  ����fU  gYL��  ��q/       consectetur @���fU  ����fU  @��cillum dolore eu fugiat nulla pariatur ��fU  @���fU  ����fU  QCL��  2�q/       exercitation ��fU  ���fU  � �Duis aute irure dolor in rehendert in volupate velit esse U  TCL��  2�q/       exercitation ���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  VCL��  2�q/       exercitation ��fU  ���fU  0�Duis aute irure dolor in rehendert in volupate velit esse U  XCL��  2�q/       exercitation I��fU  �J��fU  @K�Duis aute irure dolor in rehendert in volupate velit esse U  .�!L��  ��q/      Workout     p���fU  0���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  p��fU  0��fU  ���L��  ��q/      Meeting                        Excepteur sint occaecat cupidatat non proident               (a�L��  ��q/       consectetur                    ullamco laboris nisi ut aliquip ex ea commodo consequat      +a�L��  ��q/       consectetur �y��fU   z��fU  �z�ullamco laboris nisi ut aliquip ex ea commodo consequat e U  -a�L��  ��q/       consectetur ����fU  ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat e U  /a�L��  ��q/       consectetur ���fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat e U  ���L��  b�q/       malorum fU  P���fU  ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ���L��  b�q/       malorum ent `���fU   ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ���L��  b�q/       malorum ent 0���fU  ����fU  0��Duis aute irure dolor in rehendert in volupate velit esse U  ���L��  b�q/       malorum ent 0���fU  ����fU  p��Duis aute irure dolor in rehendert in volupate velit esse U  <JM��  w�q/      Birthday nt 0K��fU  �K��fU  0L�cillum dolore eu fugiat nulla pariatur roident ��fU  �O��fU  t��M��  
#r/      exercitation ���fU  ����fU  @��sunt in culpa qui offici desunt molit aim id est laborum. U  ���M��  �%r/       Meeting     p���fU   ���fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ���M��  �%r/       Meeting     ����fU  P���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��wN��  �Kr/      malorum     ���fU  ����fU  0��Excepteur sint occaecat cupidatat non proident ��fU  О��fU  �~O��  rr/       bonorum     �O��fU  @P��fU  �P�Excepteur sint occaecat cupidatat non proident ��fU   U��fU  �~O��  rr/       bonorum     ����fU  `���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  ��O��  $sr/       bonorum     ����fU  P���fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  ��O��  $sr/       bonorum ent p���fU  0���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  ��O��  $sr/       bonorum ent `���fU   ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  ��O��  $sr/       bonorum ent ����fU  ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  ql�O��  &�r/       Workout fU  <��fU  �<��fU  �=�cillum dolore eu fugiat nulla pariatur ��fU  B��fU  pL��fU  sl�O��  &�r/       Workout ent P[��fU  \��fU  �\�cillum dolore eu fugiat nulla pariatur im id est laborum. U  ul�O��  &�r/       Workout ent 0���fU  ����fU  p��cillum dolore eu fugiat nulla pariatur im id est laborum. U  xl�O��  &�r/       Workout ent  =��fU  �=��fU  `@�cillum dolore eu fugiat nulla pariatur im id est laborum. U  ��O��  %�r/       consectetur                    Lorem ipsum dolor sit amet, consectetur adipiscing elit      ��O��  %�r/       consectetur ����fU  p���fU  0��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��O��  %�r/       consectetur  ��fU  ���fU   �Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��O��  %�r/       consectetur                    Lorem ipsum dolor sit amet, consectetur adipiscing elit      �?�O��  ��r/      malorum     �,��fU  @-��fU  �-�sunt in culpa qui offici desunt molit aim id est laborum. U  �BP��  C�r/      consectetur �2��fU  P3��fU  4�Excepteur sint occaecat cupidatat non proident velit esse U  �?�P��  Z�r/      exercitation ��fU  ��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �Q��  �s/       Workout                        cillum dolore eu fugiat nulla pariatur                       �Q��  �s/       Workout     p|��fU  0}��fU  �}�cillum dolore eu fugiat nulla pariatur ��fU  0���fU  ����fU  �Q��  �s/       Workout     ����fU  ���fU  л�cillum dolore eu fugiat nulla pariatur ��fU  п��fU  ����fU  �Q��  �s/       Workout     P���fU  ���fU  p��cillum dolore eu fugiat nulla pariatur ��fU  @���fU  ���fU  ��R��  �6s/       exercitation R��fU  pS��fU  0T�Duis aute irure dolor in rehendert in volupate velit esse U  ��R��  �6s/       exercitation ���fU  ����fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  ��R��  �6s/       exercitation ���fU  ����fU  `��Duis aute irure dolor in rehendert in volupate velit esse U  ��R��  �6s/       exercitation ���fU   ���fU  `��Duis aute irure dolor in rehendert in volupate velit esse U  �R��  d\s/      exercitation ���fU  ����fU  ���cillum dolore eu fugiat nulla pariatur ��fU  P���fU  ����fU  �$rT��  ~�s/      Workout     ����fU  ����fU  `��cillum dolore eu fugiat nulla pariatur ��fU  p���fU  0���fU  �$	U��  &�s/      Appointment B��fU  pL��fU  �C�Excepteur sint occaecat cupidatat non proident ing elit �fU  H��U��  ]t/       bonorum     ����fU  ����fU  P��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  I��U��  ]t/       bonorum     ���fU  0��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ȕHV��  �Kt/       bonorum      S��fU  �S��fU  0T�sunt in culpa qui offici desunt molit aim id est laborum. U  ɕHV��  �Kt/       bonorum     ���fU   ��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  ���V��  pt/       Meeting     �x��fU  py��fU  0}�Duis aute irure dolor in rehendert in volupate velit esse U  ���V��  pt/       Meeting  nt �m��fU  `n��fU  �n�Duis aute irure dolor in rehendert in volupate velit esse    ���V��  pt/       Meeting  nt �b��fU  c��fU  �c�Duis aute irure dolor in rehendert in volupate velit esse    ���V��  pt/       Meeting  nt �t��fU  Pu��fU  �u�Duis aute irure dolor in rehendert in volupate velit esse    �>uW��  �t/       exercitation ��fU  ��fU  `�cillum dolore eu fugiat nulla pariatur roident ��fU  p'��fU  �>uW��  �t/       exercitation ��fU  ���fU  `�cillum dolore eu fugiat nulla pariatur roident ��fU   ��fU  �>uW��  �t/       exercitation ��fU   ��fU  ��cillum dolore eu fugiat nulla pariatur roident ��fU  `��fU  �>uW��  �t/       exercitation ���fU  ���fU  p��cillum dolore eu fugiat nulla pariatur roident ��fU   ���fU  L!"���  !D/      exercitation X��fU  pY��fU  0Z�Duis aute irure dolor in rehendert in volupate velit esse    �C���  J�/       consectetur  ��fU  �!��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �C���  J�/       consectetur ����fU  `���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �C���  J�/       consectetur 0��fU  ���fU  �	�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �C���  J�/       consectetur ����fU  ����fU  P��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  i�`���  ��/       bonorum tion ��fU   ��fU  ��cillum dolore eu fugiat nulla pariatur roident ��fU  �!��fU  k�`���  ��/       bonorum tion j��fU  �j��fU  �v�cillum dolore eu fugiat nulla pariatur roident onsequat iq   m�`���  ��/       bonorum tion ���fU  p���fU  0��cillum dolore eu fugiat nulla pariatur roident onsequat iq   o�`���  ��/       bonorum tion =��fU   >��fU  �>�cillum dolore eu fugiat nulla pariatur roident onsequat iq   0����  ^�/       Meeting     ���fU  �	��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   1����  ^�/       Meeting     `��fU   ��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   2����  ^�/       Meeting     ���fU  p��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   3����  ^�/       Meeting     '��fU  �'��fU  P(�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��t���  b�/       consectetur 0���fU   ���fU  P��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  ��t���  b�/       consectetur ����fU  p���fU  0��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  ��t���  b�/       consectetur 0���fU  ����fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  ��t���  b�/       consectetur `���fU  ����fU  `��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  !����  T�/       exercitation ���fU  P���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  #����  T�/       exercitation ���fU  ����fU  `��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  %����  T�/       exercitation ���fU  `���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  (����  T�/       exercitation ���fU  ���fU  Ч�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �$����  ��/      Birthday nt p���fU  ���fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �����  \�/      Appointment �9��fU  P:��fU  �1�Duis aute irure dolor in rehendert in volupate velit esse U  �����  �/       consectetur U��fU  �U��fU  Y�Excepteur sint occaecat cupidatat non proident ��fU   g��fU  �����  �/       consectetur 0���fU  ����fU  p��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �����  �/       consectetur `���fU   ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �����  �/       consectetur ����fU  ����fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ���fU  ���  �1�/       bonorum     �L��fU  �M��fU  pN�Duis aute irure dolor in rehendert in volupate velit esse U  ���  �1�/       bonorum tur P���fU  ���fU  У�Duis aute irure dolor in rehendert in volupate velit esse U  ���  �1�/       bonorum tur 0���fU  ����fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  ���  �1�/       bonorum tur  ���fU  ����fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  ,)O���  �U�/      exercitation ���fU  ����fU  p��sunt in culpa qui offici desunt molit aim id est laborum.    �$���  z}�/      consectetur  i��fU  �i��fU   j�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  HAy���  ��/       bonorum     `��fU  �`��fU  Pa�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  LAy���  ��/       bonorum     0M��fU  �M��fU  0N�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  )����  ���/       Birthday    ���fU  н��fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   -����  ���/       Birthday    ����fU  0���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �鑆��  m��/       Meeting     P���fU  ���fU  п�cillum dolore eu fugiat nulla pariatur ��fU  ����fU  P���fU  �鑆��  m��/       Meeting tur  ���fU   ���fU  ���cillum dolore eu fugiat nulla pariatur im id est laborum. U  �M����  Ȩ�/      Workout     0���fU  ����fU  `��Duis aute irure dolor in rehendert in volupate velit esse U  �g���  Xʀ/       Meeting fU  ���fU  P��fU  �Duis aute irure dolor in rehendert in volupate velit esse U  �g���  Xʀ/       Meeting fU   ��fU  ���fU   �Duis aute irure dolor in rehendert in volupate velit esse U  �g���  Xʀ/       Meeting     �o��fU  ����fU  Pq�Duis aute irure dolor in rehendert in volupate velit esse U  �g���  Xʀ/       Meeting     ����fU  `���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  r���  �ˀ/       Birthday    `p��fU   q��fU  �q�sunt in culpa qui offici desunt molit aim id est laborum. U  u���  �ˀ/       Birthday    0H��fU  �H��fU  0I�sunt in culpa qui offici desunt molit aim id est laborum. U  x���  �ˀ/       Birthday    �E��fU  pF��fU  0G�sunt in culpa qui offici desunt molit aim id est laborum. U  {���  �ˀ/       Birthday    �E��fU  `F��fU  �F�sunt in culpa qui offici desunt molit aim id est laborum. U  �����  �ˀ/       consectetur �L��fU  �M��fU  pN�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �����  �ˀ/       consectetur  T��fU   U��fU  �U�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �����  �ˀ/       consectetur  I��fU  �J��fU  @K�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �����  �ˀ/       consectetur  g��fU  �g��fU   h�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �䢇��  O�/      malorum tion ��fU  ���fU  p�sunt in culpa qui offici desunt molit aim id est laborum.    �J����  ���/       Appointment ����fU  `���fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �J����  ���/       Appointment  "��fU  0#��fU  �#�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �J����  ���/       Appointment  ���fU  `���fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �J����  ���/       Appointment  ���fU  ����fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �|O���  ~�/      malorum ent P��fU   ��fU  P�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  4�ֈ��  "=�/      Appointment U��fU  �U��fU  Y�sunt in culpa qui offici desunt molit aim id est laborum. U  ��o���  Ed�/       Meeting     p���fU  0���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��o���  Ed�/       Meeting fU  ���fU  @��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��o���  Ed�/       Meeting     l��fU  �l��fU  m�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��o���  Ed�/       Meeting     P���fU  ���fU  У�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  \�u���  �e�/       consectetur  Q��fU  �Q��fU  U�cillum dolore eu fugiat nulla pariatur ��fU  b��fU  �b��fU  ^�u���  �e�/       consectetur  q��fU  �q��fU  `r�cillum dolore eu fugiat nulla pariatur ��fU  0v��fU  �v��fU  \q}���  �g�/      bonorum fU  �x��fU  py��fU  0}�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  T}���  v��/      Meeting     ����fU  p���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �����  ���/       Appointment P��fU  ��fU  `�Duis aute irure dolor in rehendert in volupate velit esse U  	�����  ���/       Appointment                    Duis aute irure dolor in rehendert in volupate velit esse    
�����  ���/       Appointment ����fU  `���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  �����  ���/       Appointment P��fU  ���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  $k<���  8ځ/      Appointment P���fU  ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  P���fU  !HT���  T��/       Meeting     `���fU  ���fU  `��sunt in culpa qui offici desunt molit aim id est laborum. U  "HT���  T��/       Meeting      y��fU  @_��fU  �_�sunt in culpa qui offici desunt molit aim id est laborum. U  h�ы��  q �/       Appointment p%��fU  0&��fU  �&�cillum dolore eu fugiat nulla pariatur et dolor magna aliq   i�ы��  q �/       Appointment  ���fU  ����fU   ��cillum dolore eu fugiat nulla pariatur et dolor magna aliq   j�ы��  q �/       Appointment  A��fU  @B��fU  �B�cillum dolore eu fugiat nulla pariatur et dolor magna aliq   k�ы��  q �/       Appointment  G��fU  `H��fU  �H�cillum dolore eu fugiat nulla pariatur et dolor magna aliq   ��k���  �'�/      malorum                        sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �C���  �O�/       consectetur )��fU  �)��fU  @*�Duis aute irure dolor in rehendert in volupate velit esse U  �C���  �O�/       consectetur ����fU  `���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �#���  �Q�/      exercitation ���fU  @���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �����  �x�/      malorum                        sed do eiusmo tempo incidunt ut labore et dolor magna aliq   1�׎��  �Ƃ/       Workout      E��fU  �E��fU  �F�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   2�׎��  �Ƃ/       Workout tion ���fU  ���fU  л�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   |����  ʂ/      Birthday U  ���fU  P��fU  �ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  yly���  ��/       Meeting     p(��fU  0)��fU  0*�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  zly���  ��/       Meeting     7��fU  �7��fU  @8�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ,~���  -�/      Meeting     ����fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �c����  �/       consectetur @���fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �c����  �/       consectetur �=��fU  P>��fU  ?�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ������  �>�/       bonorum                        Duis aute irure dolor in rehendert in volupate velit esse    ������  �>�/       bonorum     ��fU  ���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  ������  �>�/       bonorum     ����fU  ����fU  P��Duis aute irure dolor in rehendert in volupate velit esse U  ������  �>�/       bonorum     ���fU  P��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  �<=���  �c�/       exercitation ���fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �<=���  �c�/       exercitation ���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �<=���  �c�/       exercitation ��fU  ���fU  @�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �<=���  �c�/       exercitation ��fU  ��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ܁ϑ��  ��/       malorum     0���fU  ����fU  0��cillum dolore eu fugiat nulla pariatur ��fU  ���fU  ����fU  ߁ϑ��  ��/       malorum     ����fU  p���fU   ��cillum dolore eu fugiat nulla pariatur olupate velit esse U  ��Ց��  ���/       Workout fU  ����fU  ����fU  P��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��Ց��  ���/       Workout      9��fU  @C��fU  �:�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��Ց��  ���/       Workout     ���fU  ����fU  P��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��Ց��  ���/       Workout fU   ���fU  ����fU  0�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  Uߑ��  ��/       Birthday    ����fU  ����fU   ��Excepteur sint occaecat cupidatat non proident ��fU   ���fU  Xߑ��  ��/       Birthday    ����fU  @���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �����  ���/      Appointment � ��fU  �)��fU  p"�Excepteur sint occaecat cupidatat non proident ��fU  �'��fU  |3���  _؃/      bonorum     �R��fU  pS��fU  0T�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �����  ?��/       malorum     ����fU  `���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �����  ?��/       malorum     ���fU  p��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �����  ?��/       malorum     ���fU  0��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �����  ?��/       malorum     �"��fU  `#��fU  �#�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �ɰ���  F��/      malorum                        cillum dolore eu fugiat nulla pariatur                       �i���  ���/       bonorum     p��fU  0��fU  ��cillum dolore eu fugiat nulla pariatur ��fU  ���fU  @��fU  	�i���  ���/       bonorum     0��fU  ���fU  0�cillum dolore eu fugiat nulla pariatur ��fU  ���fU  @��fU  i����  ֎/       malorum     0���fU  ����fU  0��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  ���fU  !i����  ֎/       malorum     �1��fU   2��fU  �2�cillum dolore eu fugiat nulla pariatur ��fU  6��fU  �6��fU  ����  �֎/       Appointment ?��fU  �?��fU  �@�cillum dolore eu fugiat nulla pariatur ��fU   E��fU  �E��fU  ����  �֎/       Appointment �&��fU  p'��fU  �)�cillum dolore eu fugiat nulla pariatur ��fU   5��fU  �5��fU  ����  �֎/       Appointment ����fU  ����fU   ��cillum dolore eu fugiat nulla pariatur ��fU  @���fU   ���fU  ����  �֎/       Appointment  ���fU  ����fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU  ���fU  ������  �׎/       Workout fU  4��fU  �4��fU  P5�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ������  �׎/       Workout     ����fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ������  �׎/       Workout     ����fU  ����fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ������  �׎/       Workout     ���fU   ��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �����  �!�/      consectetur  H��fU  �H��fU  �I�Excepteur sint occaecat cupidatat non proident ��fU  �M��fU  I�����  �H�/       Meeting     �<��fU  P=��fU  �=�Excepteur sint occaecat cupidatat non proident ��fU  PB��fU  J�����  �H�/       Meeting     `;��fU  �;��fU  `<�Excepteur sint occaecat cupidatat non proident ��fU  `@��fU  -˿��  �N�/      exercitation ���fU  0���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   @�]���  (t�/       Birthday                       Lorem ipsum dolor sit amet, consectetur adipiscing elit      A�]���  (t�/       Birthday    ���fU  �	��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  B�]���  (t�/       Birthday    P���fU  ����fU  P��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  C�]���  (t�/       Birthday    p���fU  ���fU  p��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ������  ���/       Birthday U  ���fU  P��fU  �sunt in culpa qui offici desunt molit aim id est laborum. U  ������  ���/       Birthday    0���fU  ����fU  0��sunt in culpa qui offici desunt molit aim id est laborum. U  ¦����  ���/       Birthday    ����fU  P���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  æ����  ���/       Birthday    @���fU  ����fU  @��sunt in culpa qui offici desunt molit aim id est laborum. U  �ʈ���  ���/       Workout                        ullamco laboris nisi ut aliquip ex ea commodo consequat      �ʈ���  ���/       Workout     `r��fU   s��fU  �s�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �ʈ���  ���/       Workout     ����fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �ʈ���  ���/       Workout     ����fU  ����fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �����  ]�/      consectetur �&��fU  p'��fU  �)�Excepteur sint occaecat cupidatat non proident ��fU  �5��fU  �P����  ��/       bonorum ent ����fU  ����fU  @��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �P����  ��/       bonorum ent 0J��fU  �J��fU  0K�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   LM����  �W�/      Meeting fU  `���fU   ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �����  �X�/       Appointment �P��fU  `Q��fU   R�Duis aute irure dolor in rehendert in volupate velit esse U  �����  �X�/       Appointment �I��fU  �J��fU  @K�Duis aute irure dolor in rehendert in volupate velit esse U  �����  �X�/       Appointment ���fU  p��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  �����  �X�/       Appointment PM��fU   N��fU  �N�Duis aute irure dolor in rehendert in volupate velit esse U  t�����  ʆ�/      bonorum     �&��fU  p'��fU  �)�Duis aute irure dolor in rehendert in volupate velit esse U  T$���  ��/      Birthday U  p���fU  0���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU  p���fU  �h����  ��/      Meeting fU  ����fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  
(i���  �A�/       Workout     @���fU   ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  (i���  �A�/       Workout fU   ���fU  ����fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  (i���  �A�/       Workout     ���fU  Ћ��fU  Џ�Duis aute irure dolor in rehendert in volupate velit esse U  (i���  �A�/       Workout     ���fU  P��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  +i����  �G�/       consectetur p���fU  0���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  /i����  �G�/       consectetur p.��fU  0/��fU  �/�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  3i����  �G�/       consectetur 0���fU  ����fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  7i����  �G�/       consectetur ���fU  ����fU  P��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �x����  �G�/       bonorum                        Excepteur sint occaecat cupidatat non proident               �x����  �G�/       bonorum ent ����fU  p���fU  P��Excepteur sint occaecat cupidatat non proident ing elit �fU  �x����  �G�/       bonorum ent �\��fU  P]��fU  ^�Excepteur sint occaecat cupidatat non proident ing elit �fU  �x����  �G�/       bonorum ent �B��fU   C��fU  �C�Excepteur sint occaecat cupidatat non proident ing elit �fU   �����  �J�/       consectetur                    Lorem ipsum dolor sit amet, consectetur adipiscing elit      �����  �J�/       consectetur  ���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  �����  �J�/       consectetur ����fU  P ��fU  �Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  �����  �J�/       consectetur ���fU  0��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  0f ���  �p�/       consectetur ���fU  `��fU   �Duis aute irure dolor in rehendert in volupate velit esse U  1f ���  �p�/       consectetur �a��fU  0b��fU  �b�Duis aute irure dolor in rehendert in volupate velit esse U  ������  3��/      Birthday    p���fU  ���fU  p��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �^����  d��/       Meeting                        sunt in culpa qui offici desunt molit aim id est laborum.    �^����  d��/       Meeting     ����fU   ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  �^����  d��/       Meeting     p���fU  ����fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  �^����  d��/       Meeting fU  ����fU  ����fU  P��sunt in culpa qui offici desunt molit aim id est laborum. U   I5���  ���/       Birthday    `>��fU  �>��fU  `?�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   I5���  ���/       Birthday    �=��fU  P>��fU  ?�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   |�v���  �	�/      exercitation -��fU  �.��fU  �C�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  1�����  ~�/       malorum     @���fU  ����fU  s�Excepteur sint occaecat cupidatat non proident ��fU  �v��fU  2�����  ~�/       malorum     P���fU  ����fU  P��Excepteur sint occaecat cupidatat non proident ��fU  н��fU  ������  ,�/      malorum fU  `���fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   1�����  T�/       Workout     p"��fU  0#��fU  �#�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  4�����  T�/       Workout     ����fU  ����fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  7�����  T�/       Workout                        ullamco laboris nisi ut aliquip ex ea commodo consequat      :�����  T�/       Workout     ���fU  ����fU  P��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  b]����  V�/       exercitation z��fU  �{��fU  `|�Duis aute irure dolor in rehendert in volupate velit esse U  e]����  V�/       exercitation ���fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  h]����  V�/       exercitation ���fU  `���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  k]����  V�/       exercitation D��fU  �D��fU  �G�Duis aute irure dolor in rehendert in volupate velit esse U  xj����  �Z�/       Meeting fU  ����fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  {j����  �Z�/       Meeting     ����fU  p���fU  0��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ~j����  �Z�/       Meeting     ���fU  Ћ��fU  Џ�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �j����  �Z�/       Meeting      ���fU  ����fU  0��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ŗ=���  \~�/      consectetur �X��fU  pY��fU  0Z�Duis aute irure dolor in rehendert in volupate velit esse U  ��>���  �~�/       Appointment ����fU  ����fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��>���  �~�/       Appointment �O��fU  @P��fU  �P�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��>���  �~�/       Appointment ����fU  ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��>���  �~�/       Appointment ����fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  |�v���  Β/      Appointment ���fU  `���fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  �� ���  ��/      Appointment ����fU  `���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  �&y���  ��/       Meeting     �+��fU  p,��fU  �,�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �&y���  ��/       Meeting     �I��fU  �J��fU  @K�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �&y���  ��/       Meeting     ?��fU  �?��fU  P@�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �&y���  ��/       Meeting     �^��fU  _��fU  �_�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ������  �d�/       consectetur 0��fU  ���fU  �	�Excepteur sint occaecat cupidatat non proident ��fU  ���fU  ������  �d�/       consectetur ����fU  ����fU  `��Excepteur sint occaecat cupidatat non proident ��fU  `���fU  ������  �d�/       consectetur P���fU  ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  P��fU  ������  �d�/       consectetur @���fU  ����fU  p��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �tF���  ҈�/      malorum                        sunt in culpa qui offici desunt molit aim id est laborum.    ������  g��/      consectetur ����fU   ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  \����  ���/      exercitation ���fU   ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  p�����  �)�/       Birthday    @��fU   ��fU  ��Duis aute irure dolor in rehendert in volupate velit esse    q�����  �)�/       Birthday    ����fU  @���fU  ���Duis aute irure dolor in rehendert in volupate velit esse    r�����  �)�/       Birthday    @���fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse    s�����  �)�/       Birthday     Q��fU  �Q��fU  U�Duis aute irure dolor in rehendert in volupate velit esse    �8����  �u�/      consectetur p���fU  0���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  `���fU  �}���  �/      bonorum     `���fU  ���fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  uO�  �  
�/      Appointment  ��fU  ���fU  � �Duis aute irure dolor in rehendert in volupate velit esse U  ��  �  *�/       bonorum                        ullamco laboris nisi ut aliquip ex ea commodo consequat      ��  �  *�/       bonorum ent ����fU  ����fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��  �  *�/       bonorum ent �5��fU  `6��fU  �6�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��  �  *�/       bonorum ent @f��fU   g��fU  �j�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �e: �  ��/      exercitation ���fU   ���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU   ���fU  y�L �  ��/       consectetur `���fU   ���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  z�L �  ��/       consectetur ����fU  `���fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  p�� �  f<�/       Workout     �_��fU  �k��fU  �a�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  q�� �  f<�/       Workout     `?��fU  @��fU  �@�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  r�� �  f<�/       Workout     =��fU  �=��fU  `>�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  s�� �  f<�/       Workout      :��fU  �:��fU  `;�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��z �  a�/      consectetur �x��fU  py��fU  0}�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ,& �  ͌�/      malorum                        Duis aute irure dolor in rehendert in volupate velit esse    �J� �  歠/      consectetur �L��fU  @M��fU   N�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  XN� �  筠/       malorum fU  �e��fU  Pf��fU  g�cillum dolore eu fugiat nulla pariatur ��fU  �j��fU  �k��fU  YN� �  筠/       malorum     0W��fU  �W��fU  �X�cillum dolore eu fugiat nulla pariatur ��fU  �\��fU  �]��fU  ZN� �  筠/       malorum     �M��fU  N��fU  �N�cillum dolore eu fugiat nulla pariatur ��fU   R��fU  �R��fU  ]N� �  筠/       malorum     �c��fU  0d��fU  �d�cillum dolore eu fugiat nulla pariatur ��fU  �g��fU  `h��fU  }� �  ʱ�/       exercitation ���fU  `���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  }� �  ʱ�/       exercitation ���fU  ����fU  p��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  0�� �  ���/       consectetur �t��fU  �u��fU   ��cillum dolore eu fugiat nulla pariatur ��fU  �z��fU  �{��fU  1�� �  ���/       consectetur �t��fU  �u��fU   ��cillum dolore eu fugiat nulla pariatur ��fU  �z��fU  �{��fU  2�� �  ���/       consectetur  i��fU  �i��fU  `j�cillum dolore eu fugiat nulla pariatur ��fU  �m��fU  `n��fU  3�� �  ���/       consectetur 0���fU  ����fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU  ����fU  �^� �  )�/       Appointment ����fU  ����fU   ��Excepteur sint occaecat cupidatat non proident ��fU   ���fU  �^� �  )�/       Appointment ���fU  ����fU  @��Excepteur sint occaecat cupidatat non proident ��fU   ���fU  ��	 �  ��/       exercitation ���fU  ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��	 �  ��/       exercitation ���fU  ����fU  `��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��	 �  ��/       exercitation ���fU  ����fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��	 �  ��/       exercitation ���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �2	 �  ��/      exercitation l��fU  �l��fU  �m�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �r0
 �  :Z�/      Birthday U  P���fU  ���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU  P���fU  (��3 �  	�/       bonorum     ����fU  @���fU  p��cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  )��3 �  	�/       bonorum     �z��fU  �{��fU  p|�cillum dolore eu fugiat nulla pariatur ommodo consequat . U  �}4 �  ^.�/      Birthday     ���fU  ����fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU  ����fU  )=�4 �  I4�/       Meeting ent P1��fU  �1��fU  P2�sunt in culpa qui offici desunt molit aim id est laborum. U  *=�4 �  I4�/       Meeting ent ���fU  Ћ��fU  Џ�sunt in culpa qui offici desunt molit aim id est laborum. U  ���5 �  ��/       Appointment `���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ���5 �  ��/       Appointment   ��fU  �)��fU  p"�Duis aute irure dolor in rehendert in volupate velit esse U  ���5 �  ��/       Appointment  =��fU  P>��fU  ?�Duis aute irure dolor in rehendert in volupate velit esse U  ���5 �  ��/       Appointment  ��fU  �	��fU   
�Duis aute irure dolor in rehendert in volupate velit esse U  ���5 �  ���/      exercitation                   sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��b6 �  ���/       Meeting     ����fU  P���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��b6 �  ���/       Meeting     �*��fU  �+��fU  P,�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��b6 �  ���/       Meeting     � ��fU  P!��fU  �!�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��b6 �  ���/       Meeting     �B��fU  pC��fU  �C�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  <��7 �  w��/      bonorum     �&��fU  p'��fU  �)�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ʌ8 �  M�/       exercitation ���fU  ����fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ͌8 �  M�/       exercitation X��fU  `o��fU  �Y�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  Ќ8 �  M�/       exercitation [��fU  \��fU  �\�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ӌ8 �  M�/       exercitation  ��fU  � ��fU  �!�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  o!8 �  
�/       exercitation ���fU  0���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  p���fU  0���fU  o!8 �  
�/       exercitation ���fU  @���fU  p��cillum dolore eu fugiat nulla pariatur roident ��fU  0���fU  o!8 �  
�/       exercitation ���fU  `���fU   ��cillum dolore eu fugiat nulla pariatur roident ��fU  `���fU  o!8 �  
�/       exercitation ���fU  @���fU  ���cillum dolore eu fugiat nulla pariatur roident ��fU  ����fU  8�!8 �  �/       exercitation ��fU  ���fU  �	�Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  ;�!8 �  �/       exercitation                   Lorem ipsum dolor sit amet, consectetur adipiscing elit .    >�!8 �  �/       exercitation ���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  A�!8 �  �/       exercitation ���fU   ���fU  P��Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  �=�9 �  I��/      bonorum                        Lorem ipsum dolor sit amet, consectetur adipiscing elit      ��; �  �߮/      Birthday                       Lorem ipsum dolor sit amet, consectetur adipiscing elit      4��; �  ��/      Workout     p%��fU  0&��fU  �&�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU   9J< �  �-�/       Workout     0���fU   ���fU  P��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  9J< �  �-�/       Workout     Pc��fU  �c��fU  �d�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  9J< �  �-�/       Workout      d��fU  �d��fU   e�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  9J< �  �-�/       Workout fU  �2��fU   3��fU  �3�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �O< �  �.�/      bonorum     '��fU  �'��fU  P(�sunt in culpa qui offici desunt molit aim id est laborum. U  ���< �  /U�/       exercitation d��fU  `e��fU   f�sunt in culpa qui offici desunt molit aim id est laborum. U  ���< �  /U�/       exercitation ���fU  ����fU  P��sunt in culpa qui offici desunt molit aim id est laborum. U  ���< �  /U�/       exercitation ���fU  ���fU  л�sunt in culpa qui offici desunt molit aim id est laborum. U  ���< �  /U�/       exercitation e��fU  0f��fU  �f�sunt in culpa qui offici desunt molit aim id est laborum. U  �t�< �  �V�/      exercitation !��fU  P"��fU  #�cillum dolore eu fugiat nulla pariatur ��fU  '��fU  �'��fU  @��= �  h��/       bonorum fU  U��fU  �U��fU  Y�cillum dolore eu fugiat nulla pariatur ��fU  @f��fU   g��fU  A��= �  h��/       bonorum tion i��fU  j��fU  �j�cillum dolore eu fugiat nulla pariatur im id est laborum. U  B��= �  h��/       bonorum tion ���fU  ���fU  ���cillum dolore eu fugiat nulla pariatur im id est laborum. U  C��= �  h��/       bonorum tion p��fU   q��fU  �q�cillum dolore eu fugiat nulla pariatur im id est laborum. U  ��? �  ��/       Birthday    P���fU  ���fU  ���cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  ��? �  ��/       Birthday nt ���fU  �	��fU  ��cillum dolore eu fugiat nulla pariatur ommodo consequat e U  ��? �  ��/       Birthday nt `���fU  ���fU  `��cillum dolore eu fugiat nulla pariatur ommodo consequat e U  ��? �  ��/       Birthday nt @���fU  ����fU  @��cillum dolore eu fugiat nulla pariatur ommodo consequat e U  �A �  j�/       exercitation #��fU  p$��fU  �$�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �A �  j�/       exercitation ���fU  p���fU  0��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  hX�A �  щ�/       Meeting     ����fU  `���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  kX�A �  щ�/       Meeting     ����fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  nX�A �  щ�/       Meeting fU  ����fU  `���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  qX�A �  щ�/       Meeting fU  P���fU  P��fU  �1�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  A�A �  ��/       malorum     �+��fU  p,��fU  �,�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  D�A �  ��/       malorum tion                   ullamco laboris nisi ut aliquip ex ea commodo consequat e    G�A �  ��/       malorum tion ���fU  p���fU  0��ullamco laboris nisi ut aliquip ex ea commodo consequat e U  J�A �  ��/       malorum tion ���fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat e U  �q�A �  D��/       bonorum     ����fU  ����fU  ���Excepteur sint occaecat cupidatat non proident ��fU  `���fU  �q�A �  D��/       bonorum fU  �^��fU  _��fU  �_�Excepteur sint occaecat cupidatat non proident ��fU  �c��fU  �q�A �  D��/       bonorum fU  `Y��fU  �Y��fU  �Z�Excepteur sint occaecat cupidatat non proident ��fU  0^��fU  �q�A �  D��/       bonorum     `j��fU  �j��fU  �v�Excepteur sint occaecat cupidatat non proident ��fU  �o��fU  x>B �  ճ�/       consectetur                    sed do eiusmo tempo incidunt ut labore et dolor magna aliq   
x>B �  ճ�/       consectetur ����fU  `���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   x>B �  ճ�/       consectetur `>��fU  �>��fU  `?�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   x>B �  ճ�/       consectetur ���fU  Ћ��fU  Џ�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   uEB �  ���/       exercitation ���fU  ����fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  xEB �  ���/       exercitation ���fU   ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU   ���fU  T*IB �  ���/       exercitation ���fU  P���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  W*IB �  ���/       exercitation t��fU   u��fU  �u�ullamco laboris nisi ut aliquip ex ea commodo consequat iq   U�LB �  v��/      Birthday    `���fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��tC �  K�/       Meeting fU  ����fU  p���fU  P��Duis aute irure dolor in rehendert in volupate velit esse U  ��tC �  K�/       Meeting     �Y��fU  �Z��fU  P[�Duis aute irure dolor in rehendert in volupate velit esse U  ��tC �  K�/       Meeting     ����fU  @���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ��tC �  K�/       Meeting     ����fU  @���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ,#5E �  v�/      exercitation 9��fU  p:��fU   =�Excepteur sint occaecat cupidatat non proident ��fU  `I��fU  �J�o �  �Q�/      Workout     ���fU  P��fU  �Excepteur sint occaecat cupidatat non proident onsequat �fU  `^p �  �p�/       consectetur p.��fU  0/��fU  �/�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   a^p �  �p�/       consectetur ���fU  �	��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   b^p �  �p�/       consectetur ����fU  ����fU  @��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   e^p �  �p�/       consectetur ����fU  @���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �*p �  lu�/       malorum     ���fU  ����fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �*p �  lu�/       malorum     �y��fU   z��fU  �z�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ϋ3p �  �w�/      malorum ent 01��fU  �1��fU  `2�ullamco laboris nisi ut aliquip ex ea commodo consequat . U  ��Oq �  d��/       Appointment p���fU  0���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ��Oq �  d��/       Appointment ���fU  ����fU  `��Duis aute irure dolor in rehendert in volupate velit esse U  ��Oq �  d��/       Appointment ����fU  ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ��Oq �  d��/       Appointment ����fU  ����fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  ���q �  ��/       Meeting      ���fU  ����fU  p��sunt in culpa qui offici desunt molit aim id est laborum. U  ���q �  ��/       Meeting     ����fU  ����fU  `��sunt in culpa qui offici desunt molit aim id est laborum. U  ���q �  �/       malorum                        Excepteur sint occaecat cupidatat non proident               ���q �  �/       malorum     `���fU   ���fU  ���Excepteur sint occaecat cupidatat non proident onsequat �fU  ���q �  �/       malorum      R��fU  �R��fU   S�Excepteur sint occaecat cupidatat non proident onsequat �fU  ���q �  �/       malorum      h��fU  �h��fU   i�Excepteur sint occaecat cupidatat non proident onsequat �fU  �I�q �  �/      bonorum     ���fU  ����fU  p��Duis aute irure dolor in rehendert in volupate velit esse U  D+�r �  ��/      exercitation 5��fU  �5��fU  �9�Duis aute irure dolor in rehendert in volupate velit esse U  ��)s �  �9�/       Appointment �`��fU  Pa��fU  b�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��)s �  �9�/       Appointment �Y��fU  Z��fU  �Z�ullamco laboris nisi ut aliquip ex ea commodo consequat e U  ��)s �  �9�/       Appointment  W��fU  �W��fU  `X�ullamco laboris nisi ut aliquip ex ea commodo consequat e U  ��)s �  �9�/       Appointment �I��fU  @J��fU  �J�ullamco laboris nisi ut aliquip ex ea commodo consequat e U  ��/s �  S;�/      Meeting     �g��fU  `h��fU   i�Duis aute irure dolor in rehendert in volupate velit esse U  �o�s �  X_�/       Birthday     5��fU  �5��fU  �9�cillum dolore eu fugiat nulla pariatur ��fU  D��fU  �D��fU  �o�s �  X_�/       Birthday U  ���fU  P��fU   �cillum dolore eu fugiat nulla pariatur et dolor magna aliq   �o�s �  X_�/       Birthday    �L��fU  @M��fU   N�cillum dolore eu fugiat nulla pariatur et dolor magna aliq   �o�s �  X_�/       Birthday     x��fU  �x��fU  �y�cillum dolore eu fugiat nulla pariatur et dolor magna aliq   ��_t �  1��/      Appointment  ���fU  ����fU  `��sunt in culpa qui offici desunt molit aim id est laborum. U   ��t �   ��/       bonorum fU  @K��fU   L��fU  �L�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��t �   ��/       bonorum tur �:��fU  �;��fU  <�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��t �   ��/       bonorum tur `<��fU   =��fU  �=�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��t �   ��/       bonorum tur  H��fU  �H��fU  0I�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   h߄u �  1Խ/       bonorum     �	��fU  p
��fU   �cillum dolore eu fugiat nulla pariatur ��fU  p��fU  0��fU  i߄u �  1Խ/       bonorum     0���fU  ����fU  ��cillum dolore eu fugiat nulla pariatur ��fU  `���fU  ����fU  \Rv �  g��/       malorum tion b��fU  �b��fU  Pc�sunt in culpa qui offici desunt molit aim id est laborum. U  `Rv �  g��/       malorum tion ���fU   ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  �cv �  0��/       exercitation ���fU  ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �cv �  0��/       exercitation ���fU  ����fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat e    �cv �  0��/       exercitation ���fU   ��fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat e    �cv �  0��/       exercitation 5��fU  �5��fU  P6�ullamco laboris nisi ut aliquip ex ea commodo consequat e    ��v �  ���/      exercitation t��fU  �u��fU   ��cillum dolore eu fugiat nulla pariatur ��fU  �z��fU  �{��fU  ��v �  ���/       bonorum tion n��fU  �n��fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat e U  ��v �  ���/       bonorum tion ���fU  ����fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat e U  ��v �  ��/       Appointment �C��fU   D��fU  �D�Duis aute irure dolor in rehendert in volupate velit esse U  ��v �  ��/       Appointment �=��fU  P>��fU  ?�Duis aute irure dolor in rehendert in volupate velit esse U  ���v �  �"�/      Appointment ����fU  @���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �v �  U#�/       Meeting fU  @K��fU   L��fU  �L�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  	�v �  U#�/       Meeting      ���fU  ����fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  
�v �  U#�/       Meeting     ����fU  @���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �v �  U#�/       Meeting     ����fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��Ow �  �I�/      Birthday    �L��fU  �M��fU  pN�sunt in culpa qui offici desunt molit aim id est laborum. U  �Sw �  �J�/       Birthday U  �s��fU  pt��fU  0u�cillum dolore eu fugiat nulla pariatur ��fU  px��fU  0y��fU  �Sw �  �J�/       Birthday     c��fU  �c��fU  �d�cillum dolore eu fugiat nulla pariatur ��fU   i��fU  �i��fU  �Sw �  �J�/       Birthday    0V��fU  �V��fU  0W�cillum dolore eu fugiat nulla pariatur ��fU  �Z��fU  0[��fU  �Sw �  �J�/       Birthday    pl��fU  �l��fU  pm�cillum dolore eu fugiat nulla pariatur ��fU  �p��fU   q��fU  ص�w �  �q�/       Meeting      ���fU  ����fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ٵ�w �  �q�/       Meeting tion ���fU  ���fU  `��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �
�x �  䚾/       Workout ent   ��fU  �)��fU  p"�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �
�x �  䚾/       Workout ent  ���fU  ���fU  `��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   k�y �  ���/       Workout tion ���fU  ����fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   m�y �  ���/       Workout tion ?��fU   @��fU  �@�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��y �  ���/       exercitation ���fU   ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ��y �  ���/       exercitation ���fU  `���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  ��y �  ���/       exercitation ���fU   ���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  ��y �  ���/       exercitation ���fU  ����fU  `��Duis aute irure dolor in rehendert in volupate velit esse U  Y7=z �  �	�/       Birthday    Ph��fU  �h��fU  �i�sunt in culpa qui offici desunt molit aim id est laborum. U  Z7=z �  �	�/       Birthday    @���fU  ����fU  @��sunt in culpa qui offici desunt molit aim id est laborum. U  ��Dz �  z�/      malorum      6��fU  �6��fU  �7�sunt in culpa qui offici desunt molit aim id est laborum. U  ��z �  D7�/      exercitation [��fU  \��fU  �\�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��q{ �  xX�/       Appointment                    sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��q{ �  xX�/       Appointment ���fU  ����fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   q{ �  xX�/       Appointment D��fU  �D��fU  �G�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Ôq{ �  xX�/       Appointment ����fU  `���fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �^| �  邿/      malorum     �=��fU   >��fU  �>�Excepteur sint occaecat cupidatat non proident ��fU  `B��fU  Ćd~ �  ��/      exercitation                   cillum dolore eu fugiat nulla pariatur                        � �  �C�/       Workout     U��fU  �U��fU  Y�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  � �  �C�/       Workout     �9��fU  �:��fU  P;�ullamco laboris nisi ut aliquip ex ea commodo consequat . U  � �  �C�/       Workout     `���fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat . U  � �  �C�/       Workout     `���fU  ���fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat . U  Y� �  �H�/       Workout                        cillum dolore eu fugiat nulla pariatur                       [� �  �H�/       Workout     D��fU  �D��fU  �G�cillum dolore eu fugiat nulla pariatur ��fU  U��fU  �U��fU  ]� �  �H�/       Workout     ����fU  ���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU  P���fU  _� �  �H�/       Workout     ���fU  `��fU   	�cillum dolore eu fugiat nulla pariatur ��fU  ���fU  P��fU  <�� �  7l�/      Meeting     ���fU   ��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   L�Ԁ �  ���/      bonorum      	��fU  ��fU  P
�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��[(�  �T
 /      Birthday     ���fU  ����fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   i8_(�  �U
 /       Meeting     ����fU   ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  j8_(�  �U
 /       Meeting     `���fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  hl�(�  Q~
 /       malorum     �!��fU  P"��fU  #�ullamco laboris nisi ut aliquip ex ea commodo consequat iq   il�(�  Q~
 /       malorum  ur �#��fU  �$��fU  p%�ullamco laboris nisi ut aliquip ex ea commodo consequat iq   jl�(�  Q~
 /       malorum  ur @*��fU  �*��fU  �+�ullamco laboris nisi ut aliquip ex ea commodo consequat iq   ll�(�  Q~
 /       malorum  ur �3��fU  4��fU  �4�ullamco laboris nisi ut aliquip ex ea commodo consequat iq   �� )�  8
 /       Workout     ���fU  Ћ��fU  Џ�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �� )�  8
 /       Workout     @���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �D�)�  ��
 /      exercitation                   Excepteur sint occaecat cupidatat non proident               ]R�*�  k�
 /      exercitation U��fU  �U��fU  Y�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  Hz�*�  ��
 /       exercitation                   sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Kz�*�  ��
 /       exercitation ���fU  0���fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Mz�*�  ��
 /       exercitation ���fU  ����fU  @��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Oz�*�  ��
 /       exercitation ���fU  ���fU  p��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Jٽ*�  �
 /       Meeting     ����fU   ���fU  P��Duis aute irure dolor in rehendert in volupate velit esse U  Lٽ*�  �
 /       Meeting     ����fU   ���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  Nٽ*�  �
 /       Meeting     0���fU  ���fU  p��Duis aute irure dolor in rehendert in volupate velit esse U  Pٽ*�  �
 /       Meeting     ����fU  ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  z#W+�  [ /       Meeting     ����fU  ����fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   }#W+�  [ /       Meeting     0���fU  ����fU  0��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �#W+�  [ /      Appointment @���fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   F[+�  j /       malorum                        sed do eiusmo tempo incidunt ut labore et dolor magna aliq   F[+�  j /       malorum     p���fU  ���fU  p��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   c+�  j /       Workout      W��fU  �W��fU  `X�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   c+�  j /       Workout     ����fU  P���fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��{,�  Oc /      Workout tur �0��fU  `1��fU   5�Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  �+-�  $� /       consectetur D��fU  �D��fU  �G�Excepteur sint occaecat cupidatat non proident ��fU  �U��fU  �+-�  $� /       consectetur ����fU  ����fU  @��Excepteur sint occaecat cupidatat non proident ��fU  `���fU  �+-�  $� /       consectetur p���fU  0���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  0���fU  �+-�  $� /       consectetur P$��fU  �$��fU  �%�Excepteur sint occaecat cupidatat non proident ��fU  *��fU  ��0-�  �� /      malorum     �&��fU  p'��fU  �)�sunt in culpa qui offici desunt molit aim id est laborum. U  (6K.�  �� /       consectetur D��fU  �D��fU  �G�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ,6K.�  �� /       consectetur ����fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  /6K.�  �� /       consectetur ?��fU  �?��fU  �@�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  46K.�  �� /       consectetur �o��fU  �p��fU   q�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  'X.�  9� /      consectetur p���fU  0���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   R0Y.�  }� /       Meeting     ���fU  н��fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  W0Y.�  }� /       Meeting tion ���fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse    ��Y.�  �� /       Appointment ���fU   ��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  ��Y.�  �� /       Appointment D��fU  �D��fU  �G�sunt in culpa qui offici desunt molit aim id est laborum. U  Z.�  �� /       bonorum     `���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ƓZ.�  �� /       bonorum     ����fU  P���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ɓZ.�  �� /       bonorum     ���fU   ��fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ΓZ.�  �� /       bonorum     ����fU  ����fU  p��Duis aute irure dolor in rehendert in volupate velit esse U  Qp\.�  R� /       Workout     @���fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Up\.�  R� /       Workout     ���fU  ���fU  p�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Xp\.�  R� /       Workout      ��fU  ���fU  `��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ]p\.�  R� /       Workout     `���fU   ���fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ���.�  ) /      Appointment P���fU  ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  \ʁ/�  k) /      Workout                        ullamco laboris nisi ut aliquip ex ea commodo consequat      �9'0�  �S /       Appointment ���fU  Ћ��fU  Џ�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �9'0�  �S /       Appointment ����fU  ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �9'0�  �S /       Appointment �\��fU  �]��fU  p^�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �9'0�  �S /       Appointment ����fU  ����fU  0��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��0�  w /       bonorum     �R��fU  pS��fU  0T�cillum dolore eu fugiat nulla pariatur ��fU  �X��fU  pY��fU  ��0�  w /       bonorum      ���fU  ����fU  ���cillum dolore eu fugiat nulla pariatur ��fU  `���fU   ���fU  ��0�  w /       bonorum     ����fU  ����fU   ��cillum dolore eu fugiat nulla pariatur ��fU  @���fU   ���fU  ��0�  w /       bonorum     ����fU  ����fU  0"�cillum dolore eu fugiat nulla pariatur ��fU  ����fU  `���fU  ���0�  H{ /      bonorum                        Duis aute irure dolor in rehendert in volupate velit esse    ��`1�  � /       Meeting fU  @��fU   ��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  ��`1�  � /       Meeting     �}��fU  `~��fU   �Duis aute irure dolor in rehendert in volupate velit esse U  ��`1�  � /       Meeting     D��fU  �D��fU  �G�Duis aute irure dolor in rehendert in volupate velit esse U  ��`1�  � /       Meeting     �u��fU  Pv��fU  �v�Duis aute irure dolor in rehendert in volupate velit esse U  \��1�  �� /      Birthday    ���fU  p���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �*3�   /      bonorum     D��fU  �D��fU  �G�Duis aute irure dolor in rehendert in volupate velit esse U  �Ҩ3�  �9 /       Appointment @���fU  ����fU  p��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �Ҩ3�  �9 /       Appointment ����fU  ����fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �jS4�  :e /       Workout fU   ��fU  ���fU   �sunt in culpa qui offici desunt molit aim id est laborum. U  �jS4�  :e /       Workout     P��fU  ���fU  � �sunt in culpa qui offici desunt molit aim id est laborum. U  �	5�  � /       malorum     ����fU  p���fU  P��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  �	5�  � /       malorum     ���fU  `���fU  ��Excepteur sint occaecat cupidatat non proident t laborum. U  �	5�  � /       malorum      ���fU  ����fU  `��Excepteur sint occaecat cupidatat non proident t laborum. U  �	5�  � /       malorum     ����fU  ����fU  ���Excepteur sint occaecat cupidatat non proident t laborum. U  Ъ�5�  � /       Workout     ����fU  ����fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  Ӫ�5�  � /       Workout     0s��fU  �s��fU  �x�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ժ�5�  � /       Workout     p"��fU  0#��fU  �#�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ת�5�  � /       Workout     �\��fU  P]��fU  ^�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ~��5�  � /      Meeting tur �d��fU  `e��fU   f�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  g�6�  |� /       Appointment ����fU   ��fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   j�6�  |� /       Appointment P���fU  Н��fU  P��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �w6�  �� /       malorum     D��fU  �D��fU  �G�Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  �w6�  �� /       malorum ent ����fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit e    �w6�  �� /       malorum ent `���fU  ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit e    �w6�  �� /       malorum ent ���fU  ����fU  0��Lorem ipsum dolor sit amet, consectetur adipiscing elit e    ��6�  �� /       Meeting                        ullamco laboris nisi ut aliquip ex ea commodo consequat      ��6�  �� /       Meeting     P���fU  ���fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat iq   ��6�  �� /       Meeting     ���fU  ����fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat iq   ��6�  �� /       Meeting     ����fU  0���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat iq   f�!6�  �� /      consectetur  ���fU  ����fU  `��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  lG�6�  5� /      exercitation                   cillum dolore eu fugiat nulla pariatur                       Q@�6�  R  /       malorum     g��fU  �g��fU  Ph�Duis aute irure dolor in rehendert in volupate velit esse U  R@�6�  R  /       malorum tur �A��fU  @B��fU  �B�Duis aute irure dolor in rehendert in volupate velit esse U  0�W7�  �* /       Birthday U   ��fU  ���fU  � �cillum dolore eu fugiat nulla pariatur ��fU  p%��fU  0&��fU  1�W7�  �* /       Birthday    ����fU  ����fU  `��cillum dolore eu fugiat nulla pariatur olupate velit esse U  2�W7�  �* /       Birthday    `���fU  ���fU  `��cillum dolore eu fugiat nulla pariatur olupate velit esse U  3�W7�  �* /       Birthday    ����fU  ����fU  @��cillum dolore eu fugiat nulla pariatur olupate velit esse U  �]�7�  �N /      exercitation ���fU  ���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU   ���fU  ���7�  R /       malorum     U��fU  �U��fU  Y�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ���7�  R /       malorum tur У��fU  ����fU  P��Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  ���7�  R /       malorum tur ����fU  `���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  ���7�  R /       malorum tur  ���fU  ����fU  0��Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  8Gf8�  3p /       Workout     U��fU  �U��fU  Y�sunt in culpa qui offici desunt molit aim id est laborum. U  9Gf8�  3p /       Workout ent p[��fU  0\��fU  �\�sunt in culpa qui offici desunt molit aim id est laborum. U  :Gf8�  3p /       Workout ent ����fU  ����fU   ��sunt in culpa qui offici desunt molit aim id est laborum. U  ;Gf8�  3p /       Workout ent  V��fU  �V��fU   W�sunt in culpa qui offici desunt molit aim id est laborum. U   �9�  4� /       Workout      ��fU  ���fU  P�Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  !�9�  4� /       Workout     0"��fU  �"��fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit .    T<:�  v� /      exercitation ���fU  `���fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  4u�c�  "� /      Meeting     P���fU  ����fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ���fU  \7�d�  �� /      bonorum fU  P���fU  ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  e�e�  @� /      Appointment ����fU  `���fU   ��cillum dolore eu fugiat nulla pariatur ��fU   ���fU  ����fU  �=e�  �� /       consectetur 0��fU  ���fU  �	�Duis aute irure dolor in rehendert in volupate velit esse U  �=e�  �� /       consectetur P5��fU  �5��fU  P6�Duis aute irure dolor in rehendert in volupate velit esse U  �=e�  �� /       consectetur �*��fU  �+��fU  P,�Duis aute irure dolor in rehendert in volupate velit esse U  �=e�  �� /       consectetur �M��fU  PN��fU  �N�Duis aute irure dolor in rehendert in volupate velit esse U  �)�e�  s /      Appointment  ���fU  ���fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat iq   ��lf�  }8 /      Appointment  f��fU  �f��fU  �g�cillum dolore eu fugiat nulla pariatur ��fU  �v��fU  `w��fU  :�f�  W /      bonorum     p^��fU  0_��fU  �_�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ܇g�  �~ /      Meeting                        Lorem ipsum dolor sit amet, consectetur adipiscing elit      A�h�  ȥ /       Appointment ���fU  Ћ��fU  Џ�cillum dolore eu fugiat nulla pariatur ��fU  p���fU  0���fU  C�h�  ȥ /       Appointment �!��fU  P"��fU  #�cillum dolore eu fugiat nulla pariatur ��fU  '��fU  �'��fU  E�h�  ȥ /       Appointment p���fU  0���fU  ��cillum dolore eu fugiat nulla pariatur ��fU   ���fU  ���fU  G�h�  ȥ /       Appointment  ���fU  ���fU  `��cillum dolore eu fugiat nulla pariatur ��fU  `���fU  ���fU  �@h�  �� /      malorum ent                    cillum dolore eu fugiat nulla pariatur roident               �.,h�  � /       Appointment p���fU  0���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �.,h�  � /       Appointment `j��fU  �j��fU  �v�Duis aute irure dolor in rehendert in volupate velit esse U  �.,h�  � /       Appointment  e��fU  �e��fU   f�Duis aute irure dolor in rehendert in volupate velit esse U  �.,h�  � /       Appointment `���fU   ���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  �Ui�  � /       Workout     ��fU  ���fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  �Ui�  � /       Workout     ���fU  @��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  �ei�  %� /       consectetur 0s��fU  �s��fU  �x�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �ei�  %� /       consectetur  Z��fU  [��fU  �[�Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  <Ifi�  w� /      Appointment ����fU  p���fU  P��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  A��i�  � /       exercitation ���fU  P���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  C��i�  � /       exercitation ���fU  ����fU  p��sunt in culpa qui offici desunt molit aim id est laborum.    E��i�  � /       exercitation ,��fU  �-��fU  p.�sunt in culpa qui offici desunt molit aim id est laborum.    G��i�  � /       exercitation ��fU  0��fU  ��sunt in culpa qui offici desunt molit aim id est laborum.    P��i�  � /       malorum                        ullamco laboris nisi ut aliquip ex ea commodo consequat      ���i�  9! /       Workout     ����fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ���i�  9! /       Workout     �+��fU  PM��fU  �,�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ���i�  9! /       Workout     ��fU  ���fU  P�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ���i�  9! /       Workout     ��fU  ���fU  p�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �؏j�  �G /       exercitation t��fU  �t��fU  u�cillum dolore eu fugiat nulla pariatur ��fU  @x��fU  �x��fU  �؏j�  �G /       exercitation ��fU  ���fU  P�cillum dolore eu fugiat nulla pariatur ��fU  ���fU   ��fU  ��,k�  �o /      bonorum     ���fU  Ћ��fU  Џ�cillum dolore eu fugiat nulla pariatur ��fU  p���fU  0���fU  X��k�  � /       Birthday U  p���fU  ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Y��k�  � /       Birthday    ����fU  ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Z��k�  � /       Birthday    ����fU  ����fU  P��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   \��k�  � /       Birthday    ����fU  ����fU  0��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ���k�  �� /      Meeting     � ��fU   ��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  t�Hl�  �� /      consectetur �&��fU  p'��fU  �)�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �M�l�  t� /      consectetur 0���fU  ����fU  0��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  X�l�  �� /       malorum     p���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  Z�l�  �� /       malorum     ���fU  `���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �Ԏm�  � /      Workout     0
��fU  �
��fU  0�Duis aute irure dolor in rehendert in volupate velit esse U   i
n�  �+ /       bonorum     ����fU  P���fU  ��cillum dolore eu fugiat nulla pariatur ��fU  P���fU  Х��fU  i
n�  �+ /       bonorum     p���fU  0���fU  ��cillum dolore eu fugiat nulla pariatur ��fU  0���fU   ���fU  i
n�  �+ /       bonorum     ����fU  `���fU   ��cillum dolore eu fugiat nulla pariatur ��fU  P���fU  Н��fU  i
n�  �+ /       bonorum      ���fU  ����fU  P��cillum dolore eu fugiat nulla pariatur ��fU  ���fU  н��fU  E�n�  l, /      malorum     ����fU  `���fU   ��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  x#�n�  [X /       consectetur  E��fU  �E��fU  �F�sunt in culpa qui offici desunt molit aim id est laborum. U  y#�n�  [X /       consectetur ���fU  @��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  z#�n�  [X /       consectetur �_��fU  �k��fU  �a�sunt in culpa qui offici desunt molit aim id est laborum. U  {#�n�  [X /       consectetur �A��fU  `B��fU  �B�sunt in culpa qui offici desunt molit aim id est laborum. U  �Go�  �| /       malorum     ����fU  ���fU  п�Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �Go�  �| /       malorum ent ���fU  Ћ��fU  Џ�Excepteur sint occaecat cupidatat non proident velit esse U  �Go�  �| /       malorum ent b��fU  �b��fU  @f�Excepteur sint occaecat cupidatat non proident velit esse U  �Go�  �| /       malorum ent  ���fU  ����fU  ���Excepteur sint occaecat cupidatat non proident velit esse U  �&Vo�  �� /       bonorum     P��fU  ���fU  P�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �&Vo�  �� /       bonorum     @���fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��]o�  r� /      Birthday    ����fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat . U  YH�p�  '� /       bonorum fU  ��fU  ���fU  P�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ZH�p�  '� /       bonorum     ����fU  p���fU  P��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  [H�p�  '� /       bonorum     ����fU  P���fU  p��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  \H�p�  '� /       bonorum     `���fU   ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��p�  '� /      Workout     ���fU  ���fU  p�Duis aute irure dolor in rehendert in volupate velit esse U  �cq�  �� /       Workout     0��fU  ���fU  0�cillum dolore eu fugiat nulla pariatur ��fU  0
��fU  �
��fU  �cq�  �� /       Workout     �&��fU  p'��fU  �)�cillum dolore eu fugiat nulla pariatur ��fU   5��fU  �5��fU  �Zq�  � /       malorum     p���fU  0���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �Zq�  � /       malorum tur  ��fU  ���fU  `�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �Zq�  � /       malorum tur 0s��fU  �s��fU  �x�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �Zq�  � /       malorum tur ���fU  0��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �}q�  �� /      malorum     �!��fU  p"��fU  �"�Duis aute irure dolor in rehendert in volupate velit esse U  C�#q�  �� /       consectetur p���fU  0���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  P���fU  G�#q�  �� /       consectetur  k��fU  �k��fU  Pl�Excepteur sint occaecat cupidatat non proident ��fU  ����fU  +�q�  � /       bonorum     @���fU  ����fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  +�q�  � /       bonorum     �_��fU  �k��fU  �a�ullamco laboris nisi ut aliquip ex ea commodo consequat . U  �u�q�  A /       Meeting                        sunt in culpa qui offici desunt molit aim id est laborum.    �u�q�  A /       Meeting     ����fU   ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  �u�q�  A /       Meeting     @f��fU   g��fU  �j�sunt in culpa qui offici desunt molit aim id est laborum. U  �u�q�  A /       Meeting     ����fU  ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  A�hs�  h� /       malorum     �s��fU  pt��fU  0u�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  C�hs�  h� /       malorum     Pg��fU  �g��fU  Ph�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  *�is�  �� /       malorum     �{��fU  `|��fU  �|�sunt in culpa qui offici desunt molit aim id est laborum. U  ,�is�  �� /       malorum     �f��fU  `g��fU  �g�sunt in culpa qui offici desunt molit aim id est laborum. U  $�os�  8� /      Workout     ����fU  ����fU   ��Excepteur sint occaecat cupidatat non proident ��fU   ���fU  Iћ��  �( /       bonorum     0H��fU  �H��fU  0I�sunt in culpa qui offici desunt molit aim id est laborum. U  Jћ��  �( /       bonorum ent @���fU  ����fU  @��sunt in culpa qui offici desunt molit aim id est laborum.    �����  Z�( /      Workout     `j��fU  �j��fU  �v�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  x�Ƞ�  )) /       Meeting fU  P
��fU  �
��fU  ��cillum dolore eu fugiat nulla pariatur ��fU  ���fU  ��fU  y�Ƞ�  )) /       Meeting     `���fU   ���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU   ���fU  z�Ƞ�  )) /       Meeting     п��fU  ����fU  P��cillum dolore eu fugiat nulla pariatur ��fU  P���fU  ����fU  {�Ƞ�  )) /       Meeting      ���fU  ����fU   ��cillum dolore eu fugiat nulla pariatur ��fU  p���fU  ����fU  rp��  T) /       Birthday    p���fU  ����fU  p��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   	rp��  T) /       Birthday    �o��fU   p��fU  �p�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   T��  �r) /      bonorum     ����fU  `���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU   ���fU  ����  �t) /       malorum fU  p���fU  0���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ����  �t) /       malorum ent pw��fU  �w��fU  px�Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   ����  �t) /       malorum ent  ���fU  ����fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   ����  �t) /       malorum ent p���fU   ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   �#���  ,�) /       malorum     0Z��fU  �Z��fU  p[�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �#���  ,�) /       malorum tion @��fU  �@��fU  �A�Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   T	���  ��) /      Birthday U  p%��fU  0&��fU  �&�Duis aute irure dolor in rehendert in volupate velit esse U  |B4��  ��) /      Birthday    ����fU  `���fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   `���  �6* /       exercitation ���fU  `���fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  b���  �6* /       exercitation `��fU  @a��fU  �a�Duis aute irure dolor in rehendert in volupate velit esse U  d���  �6* /       exercitation c��fU  �c��fU   d�Duis aute irure dolor in rehendert in volupate velit esse U  g���  �6* /       exercitation l��fU  �l��fU  `m�Duis aute irure dolor in rehendert in volupate velit esse U  �b��  e7* /       Birthday    ����fU  ����fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �b��  e7* /       Birthday    0���fU  ����fU  0��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �b��  e7* /       Birthday    pN��fU  0O��fU  �O�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �b��  e7* /       Birthday U  ����fU  0���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �����  �;* /       Workout     �}��fU   ~��fU  �~�Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �����  �;* /       Workout     (��fU  �(��fU  )�Excepteur sint occaecat cupidatat non proident ��fU  @-��fU  ;ꖥ�  d* /       consectetur s��fU  �s��fU  t�sunt in culpa qui offici desunt molit aim id est laborum.    =ꖥ�  d* /       consectetur  ��fU  ���fU  0�sunt in culpa qui offici desunt molit aim id est laborum.    �x���  yd* /       Appointment `���fU   ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �x���  yd* /       Appointment p���fU  0���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �x���  yd* /       Appointment p���fU  0���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �x���  yd* /       Appointment `���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  h�(��  q�* /       Workout fU  p���fU  0���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  i�(��  q�* /       Workout     ����fU  �	��fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  j�(��  q�* /       Workout     �j��fU  �k��fU  l�sunt in culpa qui offici desunt molit aim id est laborum. U  k�(��  q�* /       Workout     z��fU  �z��fU  {�sunt in culpa qui offici desunt molit aim id est laborum. U  c����  ��* /       consectetur `2��fU  �2��fU  `3�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  e����  ��* /       consectetur `���fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �C���  ��* /       Workout     P���fU  ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �C���  ��* /       Workout     � ��fU  P!��fU  �!�Duis aute irure dolor in rehendert in volupate velit esse U  �C���  ��* /       Workout     ���fU  ����fU  p��Duis aute irure dolor in rehendert in volupate velit esse U  �C���  ��* /       Workout     0$��fU   %��fU  �%�Duis aute irure dolor in rehendert in volupate velit esse U  � ���  �+ /      bonorum fU  �9��fU  P:��fU  �1�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �ބ��  $+ /      malorum     �x��fU  py��fU  0}�ullamco laboris nisi ut aliquip ex ea commodo consequat . U  ����  $+ /       consectetur ����fU  ���fU  ���Excepteur sint occaecat cupidatat non proident ing elit �fU  ����  $+ /       consectetur 0���fU  ����fU  `��Excepteur sint occaecat cupidatat non proident ing elit �fU  ���  �J+ /      Meeting fU  ����fU   ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  d����   n+ /      bonorum     ����fU  `���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ���fU  `��fU  �@��  ��+ /       bonorum  ur  ���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat . U  �@��  ��+ /       bonorum  ur �X��fU  Y��fU  �Y�ullamco laboris nisi ut aliquip ex ea commodo consequat . U  �@��  ��+ /       bonorum  ur `V��fU  �V��fU  �W�ullamco laboris nisi ut aliquip ex ea commodo consequat . U  �@��  ��+ /       bonorum  ur �b��fU  c��fU  �c�ullamco laboris nisi ut aliquip ex ea commodo consequat . U  F�H��  ȗ+ /       exercitation (��fU  �(��fU  P)�Excepteur sint occaecat cupidatat non proident ��fU  �.��fU  J�H��  ȗ+ /       exercitation )��fU  �)��fU  @*�Excepteur sint occaecat cupidatat non proident ��fU  P.��fU  ��P��  ڙ+ /       consectetur `j��fU  �j��fU  �v�Excepteur sint occaecat cupidatat non proident ��fU  �o��fU  ��P��  ڙ+ /       consectetur ���fU  �	��fU  ��Excepteur sint occaecat cupidatat non proident ��fU  ��fU  ��P��  ڙ+ /       consectetur `���fU   ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  й��fU  ��P��  ڙ+ /       consectetur ����fU  `���fU   ��Excepteur sint occaecat cupidatat non proident ��fU  `���fU  �xS��  }�+ /      Birthday    p���fU  ����fU  p��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  ����  E�+ /      malorum     ����fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �ď��  v�+ /       consectetur                    ullamco laboris nisi ut aliquip ex ea commodo consequat      �ď��  v�+ /       consectetur `r��fU   s��fU  �s�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �ď��  v�+ /       consectetur @���fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �ď��  v�+ /       consectetur `���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �_��  V
, /       bonorum     ����fU  `���fU   ��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  ����fU  �_��  V
, /       bonorum tion Y��fU  �Y��fU  PZ�cillum dolore eu fugiat nulla pariatur roident ��fU   ^��fU  ���  7, /      consectetur  ���fU  ���fU  `��sunt in culpa qui offici desunt molit aim id est laborum. U   :��  �X, /       consectetur  ��fU  �!��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  ":��  �X, /       consectetur ?��fU  �?��fU  P@�sunt in culpa qui offici desunt molit aim id est laborum. U  #:��  �X, /       consectetur P5��fU  �5��fU  P6�sunt in culpa qui offici desunt molit aim id est laborum. U  %:��  �X, /       consectetur `V��fU  �V��fU  �W�sunt in culpa qui offici desunt molit aim id est laborum. U  ��B��  �Z, /      bonorum fU  �j��fU  �k��fU  l�sunt in culpa qui offici desunt molit aim id est laborum. U  4iY��  �`, /       Meeting     `���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  6iY��  �`, /       Meeting     ����fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ���  )�, /      Appointment ����fU  `���fU   ��Duis aute irure dolor in rehendert in volupate velit esse U   .s��  ��, /       Workout     @-��fU   .��fU  �0�cillum dolore eu fugiat nulla pariatur ��fU   =��fU  �=��fU  .s��  ��, /       Workout fU  �M��fU  PN��fU  �N�cillum dolore eu fugiat nulla pariatur ��fU   R��fU  �R��fU  .s��  ��, /       Workout fU  �G��fU  `H��fU  �H�cillum dolore eu fugiat nulla pariatur ��fU  �L��fU  M��fU  .s��  ��, /       Workout     pN��fU  0O��fU  �O�cillum dolore eu fugiat nulla pariatur ��fU  0T��fU  �T��fU  �i��  ��, /       exercitation ���fU  � ��fU   �Duis aute irure dolor in rehendert in volupate velit esse U  �i��  ��, /       exercitation ���fU   ���fU  P��Duis aute irure dolor in rehendert in volupate velit esse    �i��  ��, /       exercitation ���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse    �i��  ��, /       exercitation ���fU  ����fU  `��Duis aute irure dolor in rehendert in volupate velit esse    �
��  ��, /      exercitation H��fU  �H��fU  �I�sunt in culpa qui offici desunt molit aim id est laborum. U  P4H��  � - /       Birthday U  л��fU  ����fU  ��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  Q4H��  � - /       Birthday    m��fU  �m��fU  n�Excepteur sint occaecat cupidatat non proident ing elit �fU  R4H��  � - /       Birthday    Pl��fU  �l��fU  Pm�Excepteur sint occaecat cupidatat non proident ing elit �fU  T4H��  � - /       Birthday U  �;��fU   <��fU  �<�Excepteur sint occaecat cupidatat non proident ing elit �fU  �}L��  �!- /       malorum     ����fU  ����fU  0��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �}L��  �!- /       malorum      ��fU  ���fU  P�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �̰�  �B- /       exercitation X��fU  pY��fU  0Z�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �̰�  �B- /       exercitation ���fU  ����fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �̰�  �B- /       exercitation ���fU  ����fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �̰�  �B- /       exercitation ���fU   ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  P>b��  k8 /       bonorum     P1��fU  �1��fU  �2�Excepteur sint occaecat cupidatat non proident ��fU  �6��fU  Q>b��  k8 /       bonorum     �/��fU  �0��fU  �9�Excepteur sint occaecat cupidatat non proident ��fU  `5��fU  R>b��  k8 /       bonorum     `3��fU   4��fU  �4�Excepteur sint occaecat cupidatat non proident ��fU  `8��fU  S>b��  k8 /       bonorum     �<��fU   =��fU  �=�Excepteur sint occaecat cupidatat non proident ��fU   A��fU  \<���  ��8 /       consectetur �v��fU  `w��fU  �w�Excepteur sint occaecat cupidatat non proident ��fU  �{��fU  ^<���  ��8 /       consectetur ����fU  ���fU  ���Excepteur sint occaecat cupidatat non proident ing elit �fU  p����  ��8 /       Meeting fU  g��fU  �g��fU  Ph�cillum dolore eu fugiat nulla pariatur ��fU  l��fU  �l��fU  q����  ��8 /       Meeting fU   ���fU  ����fU  0��cillum dolore eu fugiat nulla pariatur ��fU  0���fU  ����fU  r����  ��8 /       Meeting     `���fU  ����fU  `��cillum dolore eu fugiat nulla pariatur ��fU  `���fU  ����fU  u����  ��8 /       Meeting     P���fU  М��fU  P��cillum dolore eu fugiat nulla pariatur ��fU  ���fU  p���fU  n���  C�8 /      consectetur �'��fU  �(��fU  )�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  7���  ¶8 /      malorum                        sunt in culpa qui offici desunt molit aim id est laborum.    �I���  k�8 /       Appointment л��fU  ����fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  �I���  k�8 /       Appointment  ,��fU  �-��fU  p.�sunt in culpa qui offici desunt molit aim id est laborum.    �I���  k�8 /       Appointment  H��fU   I��fU  �I�sunt in culpa qui offici desunt molit aim id est laborum.    �I���  k�8 /       Appointment  ��fU  p��fU  ��sunt in culpa qui offici desunt molit aim id est laborum.    �)���  o�8 /       bonorum     `���fU  ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �)���  o�8 /       bonorum fU  ����fU  ����fU  @��Excepteur sint occaecat cupidatat non proident ��fU  `���fU  _a"��  ��8 /      Appointment �}��fU  �~��fU  p�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  X�9��  ��8 /       Appointment P���fU  ����fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  Y�9��  ��8 /       Appointment ���fU  @��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  Z�9��  ��8 /       Appointment ���fU  ���fU   �sunt in culpa qui offici desunt molit aim id est laborum. U  \�9��  ��8 /       Appointment ���fU   ��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  ܺV��  �,9 /      exercitation ���fU  ����fU  0��ullamco laboris nisi ut aliquip ex ea commodo consequat iq   ����  /R9 /       Meeting     ����fU  `���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ����  /R9 /       Meeting     P���fU  ���fU  п�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ����  /R9 /       Meeting      0��fU  �0��fU  P1�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ����  /R9 /       Meeting     `3��fU   4��fU  �4�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �����  �W9 /      Workout fU  @��fU   ��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  4����  �: /      Appointment                    Excepteur sint occaecat cupidatat non proident               �[���  �: /       bonorum     ����fU  ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �[���  �: /       bonorum      ���fU  ����fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   4����  b?: /      Appointment @���fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat . U  �r���  eA: /       Appointment #��fU  �#��fU  P$�Duis aute irure dolor in rehendert in volupate velit esse U  �r���  eA: /       Appointment Pr��fU  �r��fU  Ps�Duis aute irure dolor in rehendert in volupate velit esse U  �r���  eA: /       Appointment �t��fU   u��fU  �u�Duis aute irure dolor in rehendert in volupate velit esse U  �r���  eA: /       Appointment �}��fU  `~��fU  �~�Duis aute irure dolor in rehendert in volupate velit esse U  �w��  �c: /      malorum                        cillum dolore eu fugiat nulla pariatur                       �&��  �g: /       consectetur  ���fU  ����fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �&��  �g: /       consectetur                    Lorem ipsum dolor sit amet, consectetur adipiscing elit .    fF��  ı: /      Birthday    P���fU  ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  P���fU  �>��  �*; /       Birthday    @��fU   ��fU  ��Excepteur sint occaecat cupidatat non proident ��fU  �!��fU  �>��  �*; /       Birthday    ���fU  ����fU  P��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �>��  �*; /       Birthday    Ш��fU  ����fU  ��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �>��  �*; /       Birthday U  ����fU  ����fU  @��Excepteur sint occaecat cupidatat non proident ��fU  `���fU  @����  hT; /       malorum     �1��fU  �2��fU  `3�Duis aute irure dolor in rehendert in volupate velit esse U  A����  hT; /       malorum     ���fU   ��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  D+C��  �u; /      consectetur                    Excepteur sint occaecat cupidatat non proident               acD��  �u; /       consectetur p���fU  0���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  ccD��  �u; /       consectetur ���fU   ��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  ecD��  �u; /       consectetur p���fU  ����fU  � �Duis aute irure dolor in rehendert in volupate velit esse U  gcD��  �u; /       consectetur ����fU  P���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �I��  w; /       malorum                        Lorem ipsum dolor sit amet, consectetur adipiscing elit      �I��  w; /       malorum                        Lorem ipsum dolor sit amet, consectetur adipiscing elit      �I��  w; /       malorum     ���fU  p���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �I��  w; /       malorum     @���fU  ����fU  `��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  Pl���  �< /       Workout                        sed do eiusmo tempo incidunt ut labore et dolor magna aliq   mf���  �< /      Meeting      5��fU  �5��fU  �9�cillum dolore eu fugiat nulla pariatur ��fU  D��fU  �D��fU  �`x��  P�< /      Meeting fU  ����fU  ����fU  @��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  `���fU  ���  �[G /       exercitation ���fU  ����fU  0��Excepteur sint occaecat cupidatat non proident velit esse U  ���  �[G /       exercitation ���fU  ���fU  ���Excepteur sint occaecat cupidatat non proident velit esse U  �T�  .�G /      Birthday    Ш��fU  ����fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  Y�\�  G�G /       bonorum     U��fU  �U��fU  Y�Excepteur sint occaecat cupidatat non proident ��fU   g��fU  [�\�  G�G /       bonorum ent  ���fU  0���fU  ��Excepteur sint occaecat cupidatat non proident velit esse    ]�\�  G�G /       bonorum ent  ���fU  ����fU  0��Excepteur sint occaecat cupidatat non proident velit esse    `�\�  G�G /       bonorum ent                    Excepteur sint occaecat cupidatat non proident velit esse    �m�  ��G /       Birthday    ����fU  ����fU  `��Excepteur sint occaecat cupidatat non proident ��fU  0���fU  �m�  ��G /       Birthday    P��fU  ���fU  ��Excepteur sint occaecat cupidatat non proident ��fU  �/��fU  �m�  ��G /       Birthday    ���fU  @��fU  ��Excepteur sint occaecat cupidatat non proident ��fU  p#��fU  �m�  ��G /       Birthday    ����fU  @���fU  ���Excepteur sint occaecat cupidatat non proident ��fU   ���fU  pݢ�  ��G /       Appointment 0T��fU  �T��fU  `U�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  qݢ�  ��G /       Appointment  S��fU  �S��fU  �T�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �:1�  8�G /       Workout     ���fU  P��fU  �sunt in culpa qui offici desunt molit aim id est laborum. U  �:1�  8�G /       Workout     P���fU  О��fU  P��sunt in culpa qui offici desunt molit aim id est laborum. U  L���  �H /      Meeting     @���fU   ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �ic�  �JH /      consectetur  6��fU  �6��fU  �7�Duis aute irure dolor in rehendert in volupate velit esse U  �҈�  ��H /       malorum fU  p���fU  0���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  p���fU  �҈�  ��H /       malorum ent ����fU   ���fU  ���Excepteur sint occaecat cupidatat non proident velit esse U  �҈�  ��H /       malorum ent �B��fU  PY��fU  �D�Excepteur sint occaecat cupidatat non proident velit esse U  �҈�  ��H /       malorum ent �_��fU  @`��fU  �`�Excepteur sint occaecat cupidatat non proident velit esse U  ]���  K�H /      Workout fU  P@��fU  A��fU  �A�cillum dolore eu fugiat nulla pariatur ��fU  �E��fU  �F��fU  �\'�  M�H /       exercitation ��fU  ���fU  @�ullamco laboris nisi ut aliquip ex ea commodo consequat e U  �\'�  M�H /       exercitation ���fU  ����fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat e U  +��  ��H /      Appointment ���fU  P��fU  �ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  lP�  Y
I /      Birthday    P���fU  О��fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �i^�  �I /       bonorum     ����fU  p���fU  P��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �i^�  �I /       bonorum tur ���fU  ����fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  �i^�  �I /       bonorum tur p���fU  ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  �i^�  �I /       bonorum tur ����fU  0���fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  �^��  �4I /      consectetur ����fU  ����fU  `��Duis aute irure dolor in rehendert in volupate velit esse U  (r}�  iWI /       Workout     ����fU  ����fU  `��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  )r}�  iWI /       Workout tion H��fU  �H��fU  0I�Excepteur sint occaecat cupidatat non proident t laborum. U  b�#�  ��I /       Appointment ����fU  p���fU  0��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  d�#�  ��I /       Appointment �i��fU  j��fU  �j�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  f�#�  ��I /       Appointment �7��fU  `8��fU   9�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  h�#�  ��I /       Appointment  k��fU  P��fU  0l�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �<*�  ��I /       Appointment @��fU   ��fU  ��cillum dolore eu fugiat nulla pariatur ��fU   ��fU  �!��fU  �<*�  ��I /       Appointment  ��fU  ���fU  � �cillum dolore eu fugiat nulla pariatur roident velit esse U  �<*�  ��I /       Appointment  W��fU  �W��fU  �X�cillum dolore eu fugiat nulla pariatur roident velit esse U  �<*�  ��I /       Appointment  ��fU  ���fU  0�cillum dolore eu fugiat nulla pariatur roident velit esse U  -&3�  �I /      consectetur ���fU  P��fU  �Excepteur sint occaecat cupidatat non proident ��fU  P��fU  ~��  ?�I /       Appointment  H��fU  �H��fU  �I�sunt in culpa qui offici desunt molit aim id est laborum. U  ~��  ?�I /       Appointment ���fU  ����fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  �o��  שI /       Meeting     `j��fU  �j��fU  �v�Excepteur sint occaecat cupidatat non proident ��fU  �o��fU  �o��  שI /       Meeting     ����fU  @���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  @���fU  N���  A�I /      malorum     p���fU  0���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �zQ �  :�I /      Meeting tion ���fU  P���fU  ��cillum dolore eu fugiat nulla pariatur im id est laborum. U  ��� �  =�I /      Birthday U  �n��fU  �o��fU  `p�Excepteur sint occaecat cupidatat non proident ��fU  �u��fU  K�w!�  �J /       malorum     ����fU  ����fU   ��cillum dolore eu fugiat nulla pariatur ��fU  @���fU   ���fU  M�w!�  �J /       malorum      S��fU  �S��fU  �T�cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  h݈!�  �J /       Workout     P��fU  ��fU  `�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  i݈!�  �J /       Workout tion s��fU  �s��fU  �x�Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  j݈!�  �J /       Workout tion ���fU  ����fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  l݈!�  �J /       Workout tion ��fU  ��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  �!"�  $FJ /      exercitation ���fU  ����fU  `��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  `���fU  �"�  �gJ /       Workout      ���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat iq   	�"�  �gJ /       Workout     @7��fU  �7��fU  p8�ullamco laboris nisi ut aliquip ex ea commodo consequat iq   Xd`#�  ��J /       Workout     �j��fU  @k��fU  �n�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  Yd`#�  ��J /       Workout  ion l��fU  �l��fU  m�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  Zd`#�  ��J /       Workout  ion ���fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  [d`#�  ��J /       Workout  ion ���fU  ����fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �b�#�  <�J /      Meeting     p���fU  0���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �$�  �J /      Meeting tur 0L��fU  �L��fU  0M�cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  �%�  $K /       consectetur ����fU  `���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �%�  $K /       consectetur `V��fU  �V��fU  �W�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �%�  $K /       consectetur �P��fU  PQ��fU   R�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �%�  $K /       consectetur 0Z��fU  �Z��fU  p[�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �P�%�  �-K /      Meeting      W��fU  �W��fU  `X�cillum dolore eu fugiat nulla pariatur ��fU  �\��fU  P]��fU  H�>&�  �SK /       malorum fU  ���fU  P��fU  �Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  K�>&�  �SK /       malorum ent  ��fU  �!��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  M�>&�  �SK /       malorum ent ���fU  ����fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  O�>&�  �SK /       malorum ent P��fU  ���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��H&�  CVK /       Appointment P���fU  ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��H&�  CVK /       Appointment ����fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��H&�  CVK /       Appointment ���fU  ����fU  P��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��H&�  CVK /       Appointment ����fU  @���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  e�R&�  �XK /      Workout fU  ����fU  ����fU  @��sunt in culpa qui offici desunt molit aim id est laborum. U  ��&�  C�K /       malorum     ����fU  P���fU  p��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��&�  C�K /       malorum tur ���fU  ���fU   �Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   ��&�  C�K /       malorum tur 0��fU  ���fU  0�Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   ��&�  C�K /       malorum tur  ��fU  ���fU   �Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   0�o'�  ��K /       consectetur �,��fU  �-��fU  p.�Duis aute irure dolor in rehendert in volupate velit esse U  2�o'�  ��K /       consectetur ����fU  @���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ��s'�  ͢K /       Birthday    �z��fU  `{��fU  �{�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��s'�  ͢K /       Birthday    ����fU  P���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �h(�  ��K /      bonorum     `���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  |ۦ(�  _�K /      exercitation                   cillum dolore eu fugiat nulla pariatur                       ЛrR�  ��V /       consectetur �d��fU  `e��fU   f�cillum dolore eu fugiat nulla pariatur ��fU  `j��fU  �j��fU  ћrR�  ��V /       consectetur _��fU  �_��fU  �`�cillum dolore eu fugiat nulla pariatur  adipiscing elit �fU  қrR�  ��V /       consectetur P[��fU  \��fU  �\�cillum dolore eu fugiat nulla pariatur  adipiscing elit �fU  ӛrR�  ��V /       consectetur �o��fU  ����fU  Pq�cillum dolore eu fugiat nulla pariatur  adipiscing elit �fU  �ˑS�  �V /      Birthday nt  h��fU  �h��fU   i�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  9�S�  ��V /       Appointment ���fU  ����fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   :�S�  ��V /       Appointment ���fU   ��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �pU�  xhW /       consectetur �<��fU  P=��fU  �=�cillum dolore eu fugiat nulla pariatur ��fU  �A��fU  PB��fU  �pU�  xhW /       consectetur  {��fU  �{��fU  @|�cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  �pU�  xhW /       consectetur  ���fU  P���fU   ��cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  �pU�  xhW /       consectetur  ���fU  0���fU  ���cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  ��U�  όW /       bonorum                        sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��U�  όW /       bonorum     P;��fU  �;��fU  �<�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��U�  όW /       bonorum     `���fU  ����fU  `��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��U�  όW /       bonorum     �:��fU  �;��fU  <�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �V�  ^�W /      consectetur �F��fU  `G��fU  �G�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  (��V�  ɯW /       malorum fU  p���fU  0���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  )��V�  ɯW /       malorum     �&��fU  p'��fU  �)�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  *��V�  ɯW /       malorum     p��fU  0��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  +��V�  ɯW /       malorum     �B��fU  PY��fU  �D�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��2W�  ��W /       consectetur ����fU  P���fU  ��cillum dolore eu fugiat nulla pariatur ��fU  P���fU  ���fU  ��2W�  ��W /       consectetur P���fU  Н��fU  0��cillum dolore eu fugiat nulla pariatur  adipiscing elit iq   ��2W�  ��W /       consectetur p���fU  ����fU  p��cillum dolore eu fugiat nulla pariatur  adipiscing elit iq   ��2W�  ��W /       consectetur p���fU  ���fU  ���cillum dolore eu fugiat nulla pariatur  adipiscing elit iq   `[�W�  � X /       Meeting fU  ����fU  ����fU  `��sunt in culpa qui offici desunt molit aim id est laborum. U  a[�W�  � X /       Meeting     ����fU  0���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  b[�W�  � X /       Meeting fU  p���fU  ����fU  p��sunt in culpa qui offici desunt molit aim id est laborum. U  c[�W�  � X /       Meeting     ���fU  и��fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U   ?�X�  `MX /       bonorum                        ullamco laboris nisi ut aliquip ex ea commodo consequat      ?�X�  `MX /       bonorum     p���fU  0���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat iq   ?�X�  `MX /       bonorum      N��fU  �N��fU  �O�ullamco laboris nisi ut aliquip ex ea commodo consequat iq   ?�X�  `MX /       bonorum     �:��fU   ;��fU  �;�ullamco laboris nisi ut aliquip ex ea commodo consequat iq   յ�X�  �NX /      malorum ent `���fU   ���fU  ���Excepteur sint occaecat cupidatat non proident t laborum. U  ��Z�  �X /       exercitation                   Lorem ipsum dolor sit amet, consectetur adipiscing elit      ��Z�  �X /       exercitation ���fU  `���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit .    ��Z�  �X /       exercitation B��fU  PY��fU  �D�Lorem ipsum dolor sit amet, consectetur adipiscing elit .    ��Z�  �X /       exercitation 1��fU  2��fU  �2�Lorem ipsum dolor sit amet, consectetur adipiscing elit .    �Z�  Y�X /      Meeting     �B��fU  pC��fU  �C�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �.�Z�  ��X /       bonorum     P���fU  ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �.�Z�  ��X /       bonorum     P���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �.�Z�  ��X /       bonorum     ����fU  � ��fU   �Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �.�Z�  ��X /       bonorum      ��fU  ���fU  � �Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  9[�Z�  ��X /       Birthday    �n��fU  �o��fU  `p�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ;[�Z�  ��X /       Birthday    `���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  =[�Z�  ��X /       Birthday    �0��fU  `1��fU   5�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ?[�Z�  ��X /       Birthday    ����fU  ����fU  P��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  (N[�   �X /       malorum     �x��fU  `y��fU  z�cillum dolore eu fugiat nulla pariatur ��fU  �}��fU   ~��fU  (N[�   �X /       malorum     p��fU  0��fU  ��cillum dolore eu fugiat nulla pariatur ��fU  ���fU  @��fU  ��X[�  ��X /       Workout fU  �n��fU  �o��fU  `p�cillum dolore eu fugiat nulla pariatur ��fU  �t��fU  �u��fU  ��X[�  ��X /       Workout  ur �%��fU  P&��fU  '�cillum dolore eu fugiat nulla pariatur ommodo consequat e U  ��X[�  ��X /       Workout  ur P��fU  `A��fU  ��cillum dolore eu fugiat nulla pariatur ommodo consequat e U  ��X[�  ��X /       Workout  ur �Z��fU  [��fU  �[�cillum dolore eu fugiat nulla pariatur ommodo consequat e U  �X`[�  ��X /      malorum fU  ����fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  t��[�  �Y /      Birthday U  p%��fU  0&��fU  �&�sunt in culpa qui offici desunt molit aim id est laborum. U  �!�\�  �7Y /       Meeting     ���fU  и��fU  ���Excepteur sint occaecat cupidatat non proident ��fU   ���fU  �!�\�  �7Y /       Meeting tur @f��fU   g��fU  �j�Excepteur sint occaecat cupidatat non proident ing elit . U  �!�\�  �7Y /       Meeting tur `@��fU   A��fU  D�Excepteur sint occaecat cupidatat non proident ing elit . U  �!�\�  �7Y /       Meeting tur ����fU  ����fU  `��Excepteur sint occaecat cupidatat non proident ing elit . U  ܷ�\�  �<Y /      Meeting     �&��fU  p'��fU  �)�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �Z(]�  ebY /      bonorum     �9��fU  P:��fU  �1�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �,�]�  $�Y /       bonorum      h��fU  �h��fU   i�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �,�]�  $�Y /       bonorum     ���fU  `��fU  0�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   @��]�  (�Y /       Birthday    ����fU  ����fU   ��cillum dolore eu fugiat nulla pariatur ��fU  @���fU   ���fU  A��]�  (�Y /       Birthday ion ���fU  ����fU  p��cillum dolore eu fugiat nulla pariatur im id est laborum. U  B��]�  (�Y /       Birthday ion A��fU  PB��fU  �B�cillum dolore eu fugiat nulla pariatur im id est laborum. U  D��]�  (�Y /       Birthday ion l��fU  �l��fU  �m�cillum dolore eu fugiat nulla pariatur im id est laborum. U  ��?^�  ��Y /       Meeting     `��fU   ��fU  P�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��?^�  ��Y /       Meeting      ���fU  ����fU  0��Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   ��?^�  ��Y /       Meeting     ���fU  @��fU   �Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   ��?^�  ��Y /       Meeting     ��fU  ���fU  @�Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   ��@^�  ;�Y /      consectetur ����fU  ���fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  ��^�  2�Y /      Meeting     �P��fU  `Q��fU   R�Duis aute irure dolor in rehendert in volupate velit esse U  �xx_�  ��Y /       Appointment `>��fU  �>��fU  `?�Duis aute irure dolor in rehendert in volupate velit esse U  �xx_�  ��Y /       Appointment p���fU   ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �m�_�  ��Y /      bonorum     ����fU  P���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ���fU  �ڦ`�  cGZ /       Meeting fU  ���fU  Ћ��fU  Џ�Duis aute irure dolor in rehendert in volupate velit esse U  �ڦ`�  cGZ /       Meeting     �g��fU  `h��fU   i�Duis aute irure dolor in rehendert in volupate velit esse U  �ڦ`�  cGZ /       Meeting     ����fU  `���fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  �ڦ`�  cGZ /       Meeting     p���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ���`�  %KZ /      Birthday ion ��fU  @,��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  2ظ`�  �KZ /       malorum     @���fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat e U  5ظ`�  �KZ /       malorum     P���fU  ���fU  У�ullamco laboris nisi ut aliquip ex ea commodo consequat e U  8ظ`�  �KZ /       malorum     0���fU  ����fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat e U  =ظ`�  �KZ /       malorum     ����fU  ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat e U  a5�`�  MZ /       malorum     �x��fU  py��fU  0}�Excepteur sint occaecat cupidatat non proident ��fU  Ћ��fU  d5�`�  MZ /       malorum tion ^��fU  0_��fU  �_�Excepteur sint occaecat cupidatat non proident ing elit �fU  g5�`�  MZ /       malorum tion W��fU  X��fU  �X�Excepteur sint occaecat cupidatat non proident ing elit �fU  l5�`�  MZ /       malorum tion ���fU  `���fU  ��Excepteur sint occaecat cupidatat non proident ing elit �fU  �v�`�  �NZ /       Meeting     Ш��fU  ����fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �v�`�  �NZ /       Meeting      ���fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �]a�  .vZ /      Birthday U  �L��fU  @M��fU   N�Excepteur sint occaecat cupidatat non proident ��fU  �R��fU  H��a�  ��Z /       Appointment U��fU  �U��fU  Y�cillum dolore eu fugiat nulla pariatur ��fU  @f��fU   g��fU  I��a�  ��Z /       Appointment ���fU  P��fU  �cillum dolore eu fugiat nulla pariatur et dolor magna aliq   J��a�  ��Z /       Appointment 0���fU  ����fU  0��cillum dolore eu fugiat nulla pariatur et dolor magna aliq   K��a�  ��Z /       Appointment `���fU  ����fU  `��cillum dolore eu fugiat nulla pariatur et dolor magna aliq   �_c�  ��Z /      consectetur                    Excepteur sint occaecat cupidatat non proident               1&c�  ��Z /       bonorum fU   ���fU  ����fU   x�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  2&c�  ��Z /       bonorum ent `���fU   ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  3&c�  ��Z /       bonorum ent ����fU  `���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  4&c�  ��Z /       bonorum ent  ���fU  ����fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  
J�c�  [ /       exercitation }��fU  `~��fU   �ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  J�c�  [ /       exercitation D��fU  �D��fU  �G�ullamco laboris nisi ut aliquip ex ea commodo consequat iq   J�c�  [ /       exercitation ��fU  �	��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat iq   J�c�  [ /       exercitation ���fU  ����fU  P��ullamco laboris nisi ut aliquip ex ea commodo consequat iq   %֧c�  ?[ /       malorum     �M��fU  PN��fU  �N�cillum dolore eu fugiat nulla pariatur ��fU   R��fU  �R��fU  *֧c�  ?[ /       malorum     p���fU  0���fU  ���cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  `òc�  [ /      Birthday    л��fU  ����fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  8еc�  �[ /       exercitation ���fU  ����fU  `��Excepteur sint occaecat cupidatat non proident ��fU  0���fU  =еc�  �[ /       exercitation ���fU  ����fU   x�Excepteur sint occaecat cupidatat non proident ��fU  �|��fU  Aеc�  �[ /       exercitation ���fU  ����fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  Fеc�  �[ /       exercitation 
��fU  �
��fU  0�Excepteur sint occaecat cupidatat non proident ��fU   ��fU  Ҷc�  [ /       Workout     ����fU  `���fU   ��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  Ҷc�  [ /       Workout     `���fU  ����fU  ���Excepteur sint occaecat cupidatat non proident ��fU  `���fU  Ҷc�  [ /       Workout     `s��fU   t��fU  �t�Excepteur sint occaecat cupidatat non proident ��fU   z��fU  Ҷc�  [ /       Workout     ����fU  0���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  p���fU  �V�c�  7[ /       Appointment ���fU  Ћ��fU  Џ�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �V�c�  7[ /       Appointment ����fU  ����fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �V�c�  7[ /       Appointment 0���fU  ����fU  p��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �V�c�  7[ /       Appointment `���fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Đ��  ��e /      Appointment P1��fU  �1��fU  P2�Excepteur sint occaecat cupidatat non proident ��fU  `6��fU  �����  �f /      bonorum fU  P���fU  ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  (A��  �5f /       exercitation i��fU  0j��fU  �j�sunt in culpa qui offici desunt molit aim id est laborum. U  )A��  �5f /       exercitation V��fU  �V��fU   W�sunt in culpa qui offici desunt molit aim id est laborum. U  ����  ȣf /      Meeting     �&��fU  p'��fU  �)�sunt in culpa qui offici desunt molit aim id est laborum. U  0n���  ��f /       Meeting                        Lorem ipsum dolor sit amet, consectetur adipiscing elit      2n���  ��f /       Meeting     �E��fU  �F��fU   G�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  3n���  ��f /       Meeting     ���fU  p���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  4n���  ��f /       Meeting     �F��fU  @G��fU   H�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  `G���  \�f /       malorum     ���fU  ���fU  p�Excepteur sint occaecat cupidatat non proident ��fU   ��fU  aG���  \�f /       malorum     ���fU  ����fU  P��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  bG���  \�f /       malorum     P
��fU  �
��fU  ��Excepteur sint occaecat cupidatat non proident ��fU  ��fU  cG���  \�f /       malorum     �+��fU  p,��fU  �,�Excepteur sint occaecat cupidatat non proident ��fU  P:��fU  ?y���  wg /      Meeting ent �5��fU  `6��fU  �6�Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   hɒ�  �g /       Appointment ���fU  P��fU  �Duis aute irure dolor in rehendert in volupate velit esse    iɒ�  �g /       Appointment P���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse    jɒ�  �g /       Appointment `���fU  ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse    lɒ�  �g /       Appointment �0��fU  `1��fU   5�Duis aute irure dolor in rehendert in volupate velit esse    @Y��  Hhg /       bonorum                        sed do eiusmo tempo incidunt ut labore et dolor magna aliq   AY��  Hhg /       bonorum tion ��fU  ���fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   BY��  Hhg /       bonorum tion n��fU   o��fU  �o�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   DY��  Hhg /       bonorum tion ��fU  0��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   _���  �kg /      bonorum     ��fU  ���fU  p�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �$���  x�g /       malorum     ����fU   ���fU  P��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �$���  x�g /       malorum     �"��fU  p#��fU  �#�ullamco laboris nisi ut aliquip ex ea commodo consequat e U  �$���  x�g /       malorum     ���fU  ���fU  �ullamco laboris nisi ut aliquip ex ea commodo consequat e U  �$���  x�g /       malorum     ����fU  P���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat e U  �ѕ�  ��g /      Appointment ����fU  `���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ��\��  Xh /       consectetur P$��fU  �$��fU  �%�Duis aute irure dolor in rehendert in volupate velit esse U  ��\��  Xh /       consectetur `���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ¯\��  Xh /       consectetur  ���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  į\��  Xh /       consectetur 0��fU  ���fU  0�Duis aute irure dolor in rehendert in volupate velit esse U  ��e��  �	h /      Workout     p��fU  ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �~���  ;/h /      Workout     ����fU  ����fU  `��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �!z��  kPh /       malorum     0T��fU  �T��fU  pU�sunt in culpa qui offici desunt molit aim id est laborum. U  �!z��  kPh /       malorum     ���fU  ����fU   ��sunt in culpa qui offici desunt molit aim id est laborum. U  �!z��  kPh /       malorum     ���fU  Ћ��fU  Џ�sunt in culpa qui offici desunt molit aim id est laborum. U  �!z��  kPh /       malorum     ����fU  @���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  ٴ���  �Vh /       consectetur ����fU   ���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU  `���fU  ۴���  �Vh /       consectetur �7��fU  `8��fU   9�cillum dolore eu fugiat nulla pariatur et dolor magna aliq   ݴ���  �Vh /       consectetur  S��fU  �S��fU  �T�cillum dolore eu fugiat nulla pariatur et dolor magna aliq   ߴ���  �Vh /       consectetur P��fU  ���fU  P�cillum dolore eu fugiat nulla pariatur et dolor magna aliq   ���  Mwh /       bonorum                        Lorem ipsum dolor sit amet, consectetur adipiscing elit      ���  Mwh /       bonorum     '��fU  �'��fU  P(�Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  ���  Mwh /       bonorum     0���fU  ����fU  0��Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  ���  Mwh /       bonorum     �#��fU  �$��fU  p%�Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  ����  �zh /      Birthday U  @���fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  Q����  ��h /       Birthday    p%��fU  0&��fU  �&�Duis aute irure dolor in rehendert in volupate velit esse U  T����  ��h /       Birthday    ����fU   ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  W����  ��h /       Birthday                       Duis aute irure dolor in rehendert in volupate velit esse    Z����  ��h /       Birthday    ���fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  p
Ș�  �h /       Meeting     @��fU   ��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   s
Ș�  �h /       Meeting     ���fU  P��fU  �sed do eiusmo tempo incidunt ut labore et dolor magna aliq   v
Ș�  �h /       Meeting fU  � ��fU   ��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   y
Ș�  �h /       Meeting     0J��fU  �J��fU  0K�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ro̘�  �h /       bonorum fU  �j��fU  �k��fU  l�cillum dolore eu fugiat nulla pariatur ��fU  ����fU  ���fU  uo̘�  �h /       bonorum     �a��fU  pb��fU   c�cillum dolore eu fugiat nulla pariatur ��fU   f��fU  �f��fU  xo̘�  �h /       bonorum     b��fU  �b��fU  Pc�cillum dolore eu fugiat nulla pariatur ��fU  g��fU  �g��fU  {o̘�  �h /       bonorum     0T��fU  �T��fU  pU�cillum dolore eu fugiat nulla pariatur ��fU  0Z��fU  �Z��fU  �ߙ�  v�h /       Birthday    Ч��fU  P���fU  Ш�Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �ߙ�  v�h /       Birthday    ���fU  P��fU  ��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  ��ߙ�  v�h /       Birthday    ����fU  @���fU  p��Excepteur sint occaecat cupidatat non proident ��fU  0���fU  ��ߙ�  v�h /       Birthday    ���fU   ��fU  ��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  ��  `�h /       Appointment �R��fU  pS��fU  0T�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��  `�h /       Appointment ����fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat iq   ��  `�h /       Appointment ���fU  н��fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat iq   ��  `�h /       Appointment ���fU  �	��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat iq   ��u��  �i /       Appointment P���fU  ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��u��  �i /       Appointment  ��fU  ��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��u��  �i /       Appointment  ��fU  ���fU   �sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��u��  �i /       Appointment  ��fU  0��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ,*��  Bi /      Meeting tur Pr��fU  �r��fU  Ps�Duis aute irure dolor in rehendert in volupate velit esse U  }r���  �ei /      bonorum     D��fU  �D��fU  �G�Duis aute irure dolor in rehendert in volupate velit esse U  Hɺ��  gi /       Appointment ����fU  p���fU  P��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Jɺ��  gi /       Appointment P���fU  ����fU  P��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Kɺ��  gi /       Appointment ����fU  p���fU  P��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Lɺ��  gi /       Appointment ����fU  @���fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   )3C��  	�i /       Birthday nt ����fU  ����fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ,3C��  	�i /       Birthday nt p^��fU  0_��fU  �_�ullamco laboris nisi ut aliquip ex ea commodo consequat e U  .3C��  	�i /       Birthday nt 0v��fU  �v��fU  pw�ullamco laboris nisi ut aliquip ex ea commodo consequat e U  03C��  	�i /       Birthday nt �4��fU  p5��fU  �5�ullamco laboris nisi ut aliquip ex ea commodo consequat e U   �\��  ��i /       bonorum     �x��fU  py��fU  0}�sunt in culpa qui offici desunt molit aim id est laborum. U  #�\��  ��i /       bonorum     �0��fU  `1��fU   5�sunt in culpa qui offici desunt molit aim id est laborum. U  %�\��  ��i /       bonorum     ���fU  ����fU   ��sunt in culpa qui offici desunt molit aim id est laborum. U  '�\��  ��i /       bonorum     ����fU  0���fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  �7]��  ��i /      Meeting     p%��fU  0&��fU  �&�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  t���  j�i /      consectetur @f��fU   g��fU  �j�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   9ox��  3�i /       Appointment �o��fU  �p��fU   q�cillum dolore eu fugiat nulla pariatur ��fU  0u��fU  �u��fU  :ox��  3�i /       Appointment 0J��fU  �J��fU  0K�cillum dolore eu fugiat nulla pariatur ��fU  �M��fU  PN��fU  ތ��  n�i /      Birthday    ���fU  P��fU  �ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  M��  A�i /      bonorum     ���fU  ����fU  `��sed do eiusmo tempo incidunt ut labore et dolor magna aliq    ���  tj /       malorum     �t��fU  �u��fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  "���  tj /       malorum      ���fU  ����fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  1�B��  ~Nj /       Birthday U  � ��fU  p��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat . U  2�B��  ~Nj /       Birthday     ���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat . U  �E��  EOj /      Meeting      ���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ����  �wj /       consectetur ����fU  `���fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit iq    ��  �wj /       consectetur � ��fU  P��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   à��  �wj /       consectetur ����fU  ����fU  0��Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   Ġ��  �wj /       consectetur `���fU   ���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   �.��  �yj /      Meeting fU  �X��fU  pY��fU  0Z�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �X���  �"u /      Appointment P��fU  ��fU  `�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  _0��  �Ku /       Meeting     ����fU  `���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ���fU   ��fU  _0��  �Ku /       Meeting     ���fU  @��fU  ��cillum dolore eu fugiat nulla pariatur et dolor magna aliq   Q�;��  �Nu /       exercitation 4��fU   5��fU  �5�sunt in culpa qui offici desunt molit aim id est laborum. U  S�;��  �Nu /       exercitation ���fU  `���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  ҽ��  pu /       Workout     0W��fU  �W��fU  0X�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  	ҽ��  pu /       Workout     �D��fU  PE��fU   F�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  -3���  �u /      consectetur ���fU  P��fU  �Excepteur sint occaecat cupidatat non proident ��fU  ��fU  (���  ��u /       exercitation ���fU  `���fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  *���  ��u /       exercitation g��fU  `h��fU   i�sunt in culpa qui offici desunt molit aim id est laborum. U  +���  ��u /       exercitation ��fU  �	��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  ,���  ��u /       exercitation a��fU  0b��fU  �b�sunt in culpa qui offici desunt molit aim id est laborum. U  �:���  :�u /      Birthday    D��fU  �D��fU  �G�sunt in culpa qui offici desunt molit aim id est laborum. U  ��"��  v /       Meeting     �X��fU  Y��fU  �Y�cillum dolore eu fugiat nulla pariatur ��fU  �\��fU  ]��fU  ��"��  v /       Meeting     ����fU  ����fU  @��cillum dolore eu fugiat nulla pariatur ��fU  @���fU  ����fU  H����  �5v /       Meeting fU  ����fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  I����  �5v /       Meeting fU  @���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  J����  �5v /       Meeting     @f��fU   g��fU  �j�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  K����  �5v /       Meeting      ���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  e�U��  �[v /      Appointment �L��fU  �M��fU  pN�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   h�c��  1_v /       Meeting     ����fU  P���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  j�c��  1_v /       Meeting     ����fU  P���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  k�c��  1_v /       Meeting     P���fU  ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  l�c��  1_v /       Meeting     p���fU  ���fU  p��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  D:���  �v /      Appointment ����fU  @���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ����  1�v /      exercitation ���fU  `���fU   ��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  `���fU  pAN��  Fw /       consectetur ����fU  `���fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  qAN��  Fw /       consectetur ���fU   ��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  D����  ,Kw /      Appointment ����fU  ����fU  `��cillum dolore eu fugiat nulla pariatur ��fU  p���fU  0���fU  �w���  -mw /       exercitation                   cillum dolore eu fugiat nulla pariatur                       �	���  �nw /      exercitation                   sunt in culpa qui offici desunt molit aim id est laborum.    	(��  ��w /       Workout     ����fU  0���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  
(��  ��w /       Workout     ���fU   ��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  �c.��  0�w /      Meeting     ����fU  p���fU  P��cillum dolore eu fugiat nulla pariatur ��fU  P���fU  ���fU  f���  C�w /      Birthday U  @���fU   ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  Y���  '�w /       Birthday    ����fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  Z���  '�w /       Birthday    ���fU  p���fU  0��Duis aute irure dolor in rehendert in volupate velit esse U  �����  �x /       Workout     Pq��fU  �q��fU  Pr�cillum dolore eu fugiat nulla pariatur ��fU  �u��fU  0v��fU  �����  �x /       Workout  nt ^��fU  �^��fU  _�cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  ,�|��  M0x /      malorum     ���fU  p���fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �2���  �5x /       malorum     @���fU  ����fU  @��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �2���  �5x /       malorum     Pa��fU  �a��fU  �b�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   X?1��  �^x /       Birthday     ��fU  ���fU  � �Duis aute irure dolor in rehendert in volupate velit esse U  Y?1��  �^x /       Birthday    @���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  Z?1��  �^x /       Birthday    ��fU  ���fU  P�Duis aute irure dolor in rehendert in volupate velit esse U  [?1��  �^x /       Birthday    �:��fU  �;��fU  <�Duis aute irure dolor in rehendert in volupate velit esse U  t{���  �|x /      Meeting fU  ����fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �����  �|x /       bonorum     �t��fU   u��fU  �u�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �����  �|x /       bonorum      ��fU  ���fU  P�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��>��  ��x /       consectetur `��fU  ���fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  ��>��  ��x /       consectetur  *��fU  �+��fU  P,�sunt in culpa qui offici desunt molit aim id est laborum. U  ��>��  ��x /       consectetur  ���fU  ����fU  P��sunt in culpa qui offici desunt molit aim id est laborum. U  ��>��  ��x /       consectetur  -��fU  p.��fU   /�sunt in culpa qui offici desunt molit aim id est laborum. U  �VT��  �x /       exercitation +��fU  p,��fU  �,�Excepteur sint occaecat cupidatat non proident onsequat �fU  �VT��  �x /       exercitation ���fU  @���fU  ���Excepteur sint occaecat cupidatat non proident onsequat .    �VT��  �x /       exercitation ���fU  ����fU  P��Excepteur sint occaecat cupidatat non proident onsequat .    �VT��  �x /       exercitation ���fU  ���fU  л�Excepteur sint occaecat cupidatat non proident onsequat .    �����  Y�x /       exercitation @��fU  A��fU  �A�Duis aute irure dolor in rehendert in volupate velit esse U  �����  Y�x /       exercitation ?��fU  �?��fU  P@�Duis aute irure dolor in rehendert in volupate velit esse U  �����  Y�x /       exercitation ��fU  ���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  �����  Y�x /       exercitation @��fU  �@��fU  �A�Duis aute irure dolor in rehendert in volupate velit esse U  <� ��  �y /      exercitation                   sunt in culpa qui offici desunt molit aim id est laborum.    I�(��  � y /       Meeting     ���fU  p��fU  ��Excepteur sint occaecat cupidatat non proident ��fU   ��fU  J�(��  � y /       Meeting     0$��fU   %��fU  �%�Excepteur sint occaecat cupidatat non proident ��fU  �)��fU  �̥��  �@y /       Birthday     5��fU  �5��fU  �9�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �̥��  �@y /       Birthday    ���fU  p���fU  0��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �̥��  �@y /       Birthday    �v��fU  `w��fU   l�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �̥��  �@y /       Birthday U  ����fU  P���fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��;��  kgy /       bonorum     0���fU  ����fU  p��Duis aute irure dolor in rehendert in volupate velit esse U  ��;��  kgy /       bonorum      ���fU  ����fU  `��Duis aute irure dolor in rehendert in volupate velit esse U  ��;��  kgy /       bonorum      ��fU  ���fU  `��Duis aute irure dolor in rehendert in volupate velit esse U  ��;��  kgy /       bonorum     ���fU  ����fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  �����  D�y /       exercitation ���fU  0���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �����  D�y /       exercitation #��fU  �#��fU  �$�Duis aute irure dolor in rehendert in volupate velit esse U  �����  N�y /       Meeting                        cillum dolore eu fugiat nulla pariatur                       �����  N�y /       Meeting     ����fU  0���fU  ���cillum dolore eu fugiat nulla pariatur et dolor magna aliq   ڀ���  w�y /       Appointment �2��fU  P3��fU  4�Duis aute irure dolor in rehendert in volupate velit esse U  ހ���  w�y /       Appointment `2��fU  �2��fU  `3�Duis aute irure dolor in rehendert in volupate velit esse U  �4���  (�y /      consectetur                    sunt in culpa qui offici desunt molit aim id est laborum.    ّ���  �y /       exercitation ��fU  @��fU   �Excepteur sint occaecat cupidatat non proident ��fU  ���fU  ݑ���  �y /       exercitation ���fU  @���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  t�m�  ʷ� /      Workout                        ullamco laboris nisi ut aliquip ex ea commodo consequat      ����  �ۄ /      Meeting     P���fU  ���fU  У�cillum dolore eu fugiat nulla pariatur ��fU  Ч��fU  P���fU  4���  b� /      bonorum      ��fU  ���fU  � �cillum dolore eu fugiat nulla pariatur ��fU  p%��fU  0&��fU  ����  �S� /      exercitation ���fU   ���fU  `��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  ��`	�  y� /       Meeting fU  P[��fU  \��fU  �\�sunt in culpa qui offici desunt molit aim id est laborum. U  ��`	�  y� /       Meeting     �F��fU  @G��fU   H�sunt in culpa qui offici desunt molit aim id est laborum. U  ��`	�  y� /       Meeting     �D��fU  `E��fU  �E�sunt in culpa qui offici desunt molit aim id est laborum. U  ��`	�  y� /       Meeting     `S��fU  0T��fU  �T�sunt in culpa qui offici desunt molit aim id est laborum. U  ��e	�  Pz� /       malorum                        Duis aute irure dolor in rehendert in volupate velit esse    ��e	�  Pz� /       malorum     �&��fU  p'��fU  �)�Duis aute irure dolor in rehendert in volupate velit esse U  ��e	�  Pz� /       malorum     P��fU  ���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  ��e	�  Pz� /       malorum     ���fU  @��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  @ g	�  �z� /       consectetur                    Lorem ipsum dolor sit amet, consectetur adipiscing elit      C g	�  �z� /       consectetur �I��fU  �J��fU  @K�Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   F g	�  �z� /       consectetur 0Z��fU  �Z��fU  p[�Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   I g	�  �z� /       consectetur �b��fU  c��fU  �c�Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   �-
�  ��� /      consectetur  ��fU  �!��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  t��
�  �ƅ /      Appointment p%��fU  0&��fU  �&�cillum dolore eu fugiat nulla pariatur ��fU  �+��fU  p,��fU  ����  �� /       Workout     ��fU  ���fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  ����  �� /       Workout     ���fU  ���fU   �sunt in culpa qui offici desunt molit aim id est laborum. U  O�K�  =8� /       Appointment P(��fU  �(��fU  P)�Duis aute irure dolor in rehendert in volupate velit esse U  R�K�  =8� /       Appointment  0��fU  �0��fU  P1�Duis aute irure dolor in rehendert in volupate velit esse U  9cQ�  �9� /       Appointment p���fU  0���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU  `���fU  ;cQ�  �9� /       Appointment `���fU   ���fU  ��cillum dolore eu fugiat nulla pariatur ��fU  `���fU   ���fU  =cQ�  �9� /       Appointment ����fU  `���fU  ���cillum dolore eu fugiat nulla pariatur ��fU   ���fU  ����fU  AcQ�  �9� /       Appointment  ���fU  ����fU   ��cillum dolore eu fugiat nulla pariatur ��fU   ���fU  ���fU  ��W�  N;� /       bonorum     ����fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ��W�  N;� /       bonorum     0���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ��W�  N;� /       bonorum     �&��fU  p'��fU  �)�Duis aute irure dolor in rehendert in volupate velit esse U  ��W�  N;� /       bonorum     ����fU  p���fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  ��[�  i<� /      Workout tur p���fU  ���fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat iq   ���  ub� /       bonorum fU  ����fU  P���fU  ��cillum dolore eu fugiat nulla pariatur ��fU  P���fU  ���fU  	���  ub� /       bonorum     p���fU  ���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ���fU  ����fU  
���  ub� /       bonorum     ����fU  � ��fU   �cillum dolore eu fugiat nulla pariatur ��fU   ��fU  ���fU  ���  ub� /       bonorum     ���fU  @��fU  ��cillum dolore eu fugiat nulla pariatur ��fU  ���fU  @ ��fU  ��  ^�� /      consectetur ���fU  P��fU  �Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ���  :Ն /       consectetur P@��fU  A��fU  �A�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ���  :Ն /       consectetur 0���fU  ����fU  0��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  LG��  �׆ /      malorum     ?��fU  �?��fU  �@�Excepteur sint occaecat cupidatat non proident  magna aliq   �:��  a؆ /       consectetur p���fU  ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �:��  a؆ /       consectetur �g��fU  @h��fU  �h�Duis aute irure dolor in rehendert in volupate velit esse U  �7��  �چ /       malorum     ���fU  ����fU  ��cillum dolore eu fugiat nulla pariatur ��fU  @���fU  ����fU  �7��  �چ /       malorum     ����fU   ���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU  @���fU  W��  `L� /       Appointment ����fU  ����fU  @��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  ����fU  W��  `L� /       Appointment �&��fU  p'��fU  �)�cillum dolore eu fugiat nulla pariatur roident ��fU  �5��fU  W��  `L� /       Appointment p���fU  ����fU  p��cillum dolore eu fugiat nulla pariatur roident ��fU  P���fU  W��  `L� /       Appointment ����fU  � ��fU   �cillum dolore eu fugiat nulla pariatur roident ��fU  ���fU  䲒�  �P� /      Appointment ����fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  W��  q� /      malorum     ���fU   ��fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  (��  �r� /       Workout fU  ����fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  )��  �r� /       Workout     p|��fU  0}��fU  �}�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  *��  �r� /       Workout fU  ����fU  @���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ,��  �r� /       Workout     P���fU  Н��fU  0��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �:��  >�� /      Birthday    U��fU  �U��fU  Y�cillum dolore eu fugiat nulla pariatur ��fU  @f��fU   g��fU  ��  j� /       Meeting ent ���fU  `��fU   	�sunt in culpa qui offici desunt molit aim id est laborum. U  ��  j� /       Meeting ent ���fU  @��fU   �sunt in culpa qui offici desunt molit aim id est laborum. U  ��  j� /       Meeting ent � ��fU  `!��fU  "�sunt in culpa qui offici desunt molit aim id est laborum. U  ��  j� /       Meeting ent 0+��fU  �+��fU  0,�sunt in culpa qui offici desunt molit aim id est laborum. U  -�  �8� /       Birthday                       ullamco laboris nisi ut aliquip ex ea commodo consequat      -�  �8� /       Birthday    ����fU  ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  -�  �8� /       Birthday    `���fU  ����fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  -�  �8� /       Birthday    ����fU  ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  d%�   9� /      exercitation <��fU  �<��fU  �=�Duis aute irure dolor in rehendert in volupate velit esse U  ����  �^� /      Workout ent 0���fU  ����fU  0��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �O�  �� /       consectetur ����fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �O�  �� /       consectetur p��fU  0��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �O�  �� /       consectetur `s��fU   t��fU  �t�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �O�  �� /       consectetur ���fU  ����fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  M��  �� /      Birthday    `���fU  ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  ����  쫈 /       Workout     `���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ���  쫈 /       Workout ent  ���fU  P���fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit .    �m��  �؈ /      bonorum fU  p���fU  0���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �e�@�  �� /      Workout ent ����fU  @���fU  ���Excepteur sint occaecat cupidatat non proident t laborum. U  zgA�  �Г /      malorum                        ullamco laboris nisi ut aliquip ex ea commodo consequat      i�yA�  qՓ /       Meeting                        sunt in culpa qui offici desunt molit aim id est laborum.    j�yA�  qՓ /       Meeting ent 0���fU  ����fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  k�yA�  qՓ /       Meeting ent 0��fU  ���fU  0�sunt in culpa qui offici desunt molit aim id est laborum. U  l�yA�  qՓ /       Meeting ent ��fU  ���fU  @�sunt in culpa qui offici desunt molit aim id est laborum. U  (}B�  I�� /       malorum     p���fU  0���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   )}B�  I�� /       malorum     �7��fU  `8��fU   9�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   *}B�  I�� /       malorum     0*��fU  �*��fU  �+�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   +}B�  I�� /       malorum     �A��fU  PB��fU  �B�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   |P�B�  � /      Meeting      ��fU  ���fU  � �cillum dolore eu fugiat nulla pariatur ��fU  p%��fU  0&��fU  �ʡB�  :!� /       Meeting     ���fU  Ћ��fU  Џ�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �ʡB�  :!� /       Meeting     ����fU  P���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ���C�  �j� /      bonorum     ����fU  @���fU  ���cillum dolore eu fugiat nulla pariatur et dolor magna aliq   (WD�  )�� /       Appointment `��fU  ���fU  ��Excepteur sint occaecat cupidatat non proident ��fU  `��fU  )WD�  )�� /       Appointment  ���fU  ���fU  ���Excepteur sint occaecat cupidatat non proident ing elit e     1�D�  ��� /       bonorum      ���fU  К��fU  P��Duis aute irure dolor in rehendert in volupate velit esse U  1�D�  ��� /       bonorum      ��fU  ���fU   �Duis aute irure dolor in rehendert in volupate velit esse U  �q�E�  �� /      exercitation ��fU  @ ��fU  � �Excepteur sint occaecat cupidatat non proident ing elit �fU  ��4F�  n� /       malorum     p���fU  0���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU  `���fU  ��4F�  n� /       malorum fU  ���fU  `��fU  ��cillum dolore eu fugiat nulla pariatur ��fU   ��fU  ���fU  ��4F�  n� /       malorum     b��fU  �b��fU  Pc�cillum dolore eu fugiat nulla pariatur ��fU  g��fU  �g��fU  ��4F�  n� /       malorum     p���fU  ���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ���fU  ����fU  x�YG�  {V� /       exercitation ��fU  ���fU  �sed do eiusmo tempo incidunt ut labore et dolor magna aliq   y�YG�  {V� /       exercitation v��fU  `w��fU   l�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��H�  ã� /      Appointment @��fU   ��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �PYJ�  �� /       Workout     @���fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �PYJ�  �� /       Workout     �R��fU  pS��fU  0T�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �PYJ�  �� /       Workout     m��fU  �m��fU  n�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �PYJ�  �� /       Workout     0,��fU  �,��fU  0-�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   M�jJ�  a� /      Workout     D��fU  �D��fU  �G�cillum dolore eu fugiat nulla pariatur ��fU  U��fU  �U��fU  	�-L�  Ւ� /       exercitation ���fU  ���fU  p��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  
�-L�  Ւ� /       exercitation >��fU   ?��fU  �?�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �U/L�  I�� /      Meeting      ���fU  ����fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   l
�M�  � /      Meeting fU  D��fU  �D��fU  �G�Excepteur sint occaecat cupidatat non proident ��fU  �U��fU  ��M�  � /       Appointment �x��fU  py��fU  0}�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��M�  � /       Appointment ����fU  @���fU  p��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��M�  � /       Appointment ����fU  @���fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��M�  � /       Appointment ���fU  P��fU  �Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ���N�  �+� /      consectetur �t��fU  �u��fU   ��Excepteur sint occaecat cupidatat non proident ��fU  �{��fU  ��O�  XR� /       Meeting                        cillum dolore eu fugiat nulla pariatur                       ��O�  XR� /       Meeting ent  ���fU  ����fU   ��cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  §O�  XR� /       Meeting ent P7��fU  �7��fU  �8�cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  çO�  XR� /       Meeting ent �a��fU  `b��fU   c�cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  ą�O�  � /      Birthday nt ����fU  P���fU  Ќ�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��HP�  ��� /       Meeting     @���fU  ����fU  `��Duis aute irure dolor in rehendert in volupate velit esse U  ��HP�  ��� /       Meeting     ����fU  ����fU  0��Duis aute irure dolor in rehendert in volupate velit esse U  ��PP�  �� /       Meeting                        sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��PP�  �� /       Meeting     ����fU  ����fU  `��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��PP�  �� /       Meeting     �Z��fU  [��fU  �[�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��PP�  �� /       Meeting     ����fU  ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   4�P�  �ŗ /      Appointment ����fU  `���fU  ��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  ����fU  l�R�  5� /      consectetur ����fU  p���fU  P��Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   4R�R�  ><� /       bonorum     ����fU   ���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ���fU  ����fU  6R�R�  ><� /       bonorum     P���fU  ���fU  л�cillum dolore eu fugiat nulla pariatur ��fU  п��fU  ����fU  DA�R�  L?� /      Appointment � ��fU  �)��fU  p"�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  y��R�  ;B� /       malorum     �X��fU  pY��fU  0Z�sunt in culpa qui offici desunt molit aim id est laborum. U  z��R�  ;B� /       malorum     ���fU  ����fU  0��sunt in culpa qui offici desunt molit aim id est laborum. U  {��R�  ;B� /       malorum     `���fU  ���fU  `��sunt in culpa qui offici desunt molit aim id est laborum. U  }��R�  ;B� /       malorum     �]��fU   ^��fU  �^�sunt in culpa qui offici desunt molit aim id est laborum. U  ,l|�  �� /      malorum      f��fU  �f��fU  �g�Duis aute irure dolor in rehendert in volupate velit esse U  �}�  �� /       consectetur �O��fU  �P��fU   Q�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �}�  �� /       consectetur  ���fU  ����fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  0��}�  �>� /       bonorum fU  P���fU  ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  P���fU  1��}�  �>� /       bonorum fU  p���fU  ����fU  ���Excepteur sint occaecat cupidatat non proident ��fU  P���fU  2��}�  �>� /       bonorum      g��fU  �g��fU   h�Excepteur sint occaecat cupidatat non proident ��fU  �k��fU  3��}�  �>� /       bonorum     u��fU  �u��fU  v�Excepteur sint occaecat cupidatat non proident ��fU   z��fU  �,~�  j_� /       malorum     �i��fU  0j��fU  �j�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �,~�  j_� /       malorum     ����fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �C6~�  �a� /      exercitation ���fU  ����fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  R�C~�  Re� /       Birthday    0���fU  ����fU  0��cillum dolore eu fugiat nulla pariatur roident onsequat �fU  T�C~�  Re� /       Birthday     c��fU  �c��fU   d�cillum dolore eu fugiat nulla pariatur roident onsequat �fU   k�~�  4�� /       consectetur ����fU  `���fU  ��cillum dolore eu fugiat nulla pariatur im id est laborum. U  #k�~�  4�� /       consectetur @���fU  ����fU  ���cillum dolore eu fugiat nulla pariatur im id est laborum. U  %k�~�  4�� /       consectetur P��fU  ���fU  � �cillum dolore eu fugiat nulla pariatur im id est laborum. U  'k�~�  4�� /       consectetur <��fU  �<��fU  =�cillum dolore eu fugiat nulla pariatur im id est laborum. U  e�~�  ��� /       Meeting     p���fU  0���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   e�~�  ��� /       Meeting     P��fU  ���fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   e�~�  ��� /       Meeting     ���fU  P��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq    e�~�  ��� /       Meeting     P1��fU  �1��fU  P2�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ���~�  :�� /      Workout fU  `���fU  ����fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  ����  �ң /       Meeting  ur �C��fU  @D��fU   E�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ����  �ң /       Meeting  ur  ���fU  ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ����  �ң /       Meeting  ur @f��fU   g��fU  �j�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ����  �ң /       Meeting  ur @���fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU   C���  4�� /       exercitation ���fU  ����fU   ��cillum dolore eu fugiat nulla pariatur ��fU  @���fU   ���fU  !C���  4�� /       exercitation ���fU  ����fU  @��cillum dolore eu fugiat nulla pariatur roident ��fU  `���fU  "C���  4�� /       exercitation ���fU  ����fU   ��cillum dolore eu fugiat nulla pariatur roident ��fU  ����fU  $C���  4�� /       exercitation ���fU  К��fU  P��cillum dolore eu fugiat nulla pariatur roident ��fU  0���fU  k����  �� /       malorum     ���fU  @��fU   �ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  m����  �� /       malorum     �-��fU  p.��fU   /�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  I�0��  %� /       Workout fU  0���fU  ����fU  p��Excepteur sint occaecat cupidatat non proident ��fU  0���fU  K�0��  %� /       Workout     �9��fU  �:��fU  P;�Excepteur sint occaecat cupidatat non proident ��fU  �?��fU  M�0��  %� /       Workout fU  �+��fU  ,��fU  �,�Excepteur sint occaecat cupidatat non proident ��fU  �0��fU  P�0��  %� /       Workout      k��fU  �k��fU  Pl�Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �}7��  �&� /      Appointment �;��fU   <��fU  �<�Excepteur sint occaecat cupidatat non proident ��fU   @��fU  �>��  �(� /       exercitation                   sunt in culpa qui offici desunt molit aim id est laborum.    �>��  �(� /       exercitation ���fU  ����fU   ��sunt in culpa qui offici desunt molit aim id est laborum.    �>��  �(� /       exercitation ��fU  ���fU  `�sunt in culpa qui offici desunt molit aim id est laborum.    �>��  �(� /       exercitation ���fU  `���fU  ���sunt in culpa qui offici desunt molit aim id est laborum.    ��R��  Qo� /      malorum fU  ����fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  	%]��  �q� /       Birthday    P6��fU  �6��fU  P7�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   
%]��  �q� /       Birthday    ���fU  ����fU  @��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   p��  ��� /       exercitation ���fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  q��  ��� /       exercitation ���fU  0���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  r��  ��� /       exercitation ���fU  ����fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  s��  ��� /       exercitation ���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  }����  ߽� /      Birthday    �d��fU  `e��fU   f�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �酃�   /       consectetur ����fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  �酃�   /       consectetur ����fU  0���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �酃�   /       consectetur P���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �酃�   /       consectetur ����fU  ����fU  p��Duis aute irure dolor in rehendert in volupate velit esse U  4u���  �� /       exercitation ���fU  p���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  6u���  �� /       exercitation Z��fU  [��fU  �[�Excepteur sint occaecat cupidatat non proident ��fU  _��fU  �"��  � /       consectetur  V��fU  �V��fU   W�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �"��  � /       consectetur p���fU  0���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Ђ5��  �� /       Meeting      ��fU  ���fU   �Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ҂5��  �� /       Meeting  ion ���fU  ����fU  `��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU   nɄ�  �� /       Birthday    ����fU  p���fU  0��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  p���fU  nɄ�  �� /       Birthday U   ���fU  ����fU  P��cillum dolore eu fugiat nulla pariatur olupate velit esse U  �Dc��  "8� /       Appointment                    Excepteur sint occaecat cupidatat non proident               �Dc��  "8� /       Appointment P���fU  ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU   ���fU  �Dc��  "8� /       Appointment  ���fU  ����fU  `��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  �Dc��  "8� /       Appointment � ��fU  P��fU  ��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  �l��  �:� /      Birthday     ��fU  ���fU   �Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ����  �\� /      Appointment ����fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  bŌ��  K�� /      bonorum ent ����fU  @���fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   p���  f�� /       Meeting     @���fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  r���  f�� /       Meeting     00��fU  �0��fU  P1�ullamco laboris nisi ut aliquip ex ea commodo consequat e U  t���  f�� /       Meeting     ���fU  ����fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat e U  w���  f�� /       Meeting     ����fU  ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat e U  �蕆�  ��� /       exercitation \��fU  P]��fU  ^�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �蕆�  ��� /       exercitation ���fU  ����fU  0��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �蕆�  ��� /       exercitation ���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �蕆�  ��� /       exercitation ���fU  ����fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  t�Z��  ��� /      Birthday U  p%��fU  0&��fU  �&�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  X���  �!� /       consectetur  ���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  Y���  �!� /       consectetur ����fU  `���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  Z���  �!� /       consectetur ���fU  `���fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  \���  �!� /       consectetur ���fU  ����fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �v���  �$� /       bonorum     �*��fU   +��fU  �+�Excepteur sint occaecat cupidatat non proident ing elit �fU  �v���  �$� /       bonorum  ion ���fU  0���fU  ��Excepteur sint occaecat cupidatat non proident ing elit e U  �2w��  aC� /       bonorum     `���fU   ���fU  ���Excepteur sint occaecat cupidatat non proident ing elit �fU  �2w��  aC� /       bonorum     ����fU  ����fU  ���Excepteur sint occaecat cupidatat non proident ing elit �fU  5���  �J� /      Workout      i��fU  �i��fU   j�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   t����  j� /      Workout                        Excepteur sint occaecat cupidatat non proident               �j!��  �3� /      malorum ent �=��fU   >��fU  �>�Duis aute irure dolor in rehendert in volupate velit esse U  |DÍ�  �\� /      malorum tion "��fU  0#��fU  �#�ullamco laboris nisi ut aliquip ex ea commodo consequat iq   �����  �*� /       Birthday                       ullamco laboris nisi ut aliquip ex ea commodo consequat      �����  �*� /       Birthday U  ����fU  P���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat iq   �����  �*� /       Birthday    ����fU  `���fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat iq   �����  �*� /       Birthday    @���fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat iq   ����  W� /       consectetur @���fU   ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  ����  W� /       consectetur �O��fU  pP��fU  0Q�sunt in culpa qui offici desunt molit aim id est laborum. U  ����  W� /       consectetur P���fU  ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  ����  W� /       consectetur `���fU  ����fU  `��sunt in culpa qui offici desunt molit aim id est laborum. U  �����  �X� /      Appointment                    ullamco laboris nisi ut aliquip ex ea commodo consequat      ��7��  �|� /      consectetur p���fU  0���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  0��fU  ��չ�  P�� /      Workout                        cillum dolore eu fugiat nulla pariatur                       <#\��  �ǲ /      exercitation ���fU  ����fU  `��sunt in culpa qui offici desunt molit aim id est laborum. U  	���  �� /       Birthday    P���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  
���  �� /       Birthday    0���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �����  � /      bonorum     �x��fU  py��fU  0}�Duis aute irure dolor in rehendert in volupate velit esse U  Û��  �� /       bonorum ent  {��fU  �{��fU  @|�cillum dolore eu fugiat nulla pariatur roident ��fU  P���fU  Û��  �� /       bonorum ent  ���fU  P���fU  ���cillum dolore eu fugiat nulla pariatur roident velit esse    |Ǩ��  �� /      Meeting     ����fU  ����fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �rμ�  h� /       Birthday U  Ш��fU  ����fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �rμ�  h� /       Birthday U  �B��fU  pC��fU  �C�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �rμ�  h� /       Birthday    `���fU   ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �rμ�  h� /       Birthday    �p��fU  pq��fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  WҼ�  �h� /      exercitation ���fU  ����fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  �8c��  #�� /       malorum     ����fU  ����fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �8c��  #�� /       malorum     ����fU  �	��fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �8c��  #�� /       malorum     ����fU  ����fU  0��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �8c��  #�� /       malorum     �8��fU  �9��fU  :�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  Hg���  ݵ� /       Meeting fU  U��fU  �U��fU  Y�cillum dolore eu fugiat nulla pariatur ��fU  @f��fU   g��fU  Ig���  ݵ� /       Meeting ent  ���fU  ����fU  p��cillum dolore eu fugiat nulla pariatur ommodo consequat iq   Jg���  ݵ� /       Meeting ent  Q��fU  �Q��fU  �R�cillum dolore eu fugiat nulla pariatur ommodo consequat iq   Kg���  ݵ� /       Meeting ent  y��fU  pz��fU  �z�cillum dolore eu fugiat nulla pariatur ommodo consequat iq   DN���  lٳ /      exercitation D��fU  �D��fU  �G�Duis aute irure dolor in rehendert in volupate velit esse U  ����  �۳ /       Birthday    @���fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ����  �۳ /       Birthday U  `���fU  ����fU  `��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ����  �۳ /       Birthday    `V��fU  �V��fU  �W�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ����  �۳ /       Birthday    �b��fU  c��fU  �c�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   P+��  �� /       bonorum fU  ����fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  Q+��  �� /       bonorum      E��fU  �E��fU  �F�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  R+��  �� /       bonorum     @���fU   ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  T+��  �� /       bonorum     ����fU  @���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �J+��  �� /       Appointment ���fU  @��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat e U  �J+��  �� /       Appointment P��fU  ���fU  � �ullamco laboris nisi ut aliquip ex ea commodo consequat e U  ӿ�  �-� /       Meeting      R��fU  �R��fU   S�Excepteur sint occaecat cupidatat non proident ��fU  �V��fU  	ӿ�  �-� /       Meeting tion ���fU  ����fU   ��Excepteur sint occaecat cupidatat non proident t laborum.    =Q��  $N� /      Meeting                        Excepteur sint occaecat cupidatat non proident               `����  �z� /       malorum                        sed do eiusmo tempo incidunt ut labore et dolor magna aliq   a����  �z� /       malorum     `X��fU  `o��fU  �Y�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   b����  �z� /       malorum      f��fU  �f��fU  �g�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   c����  �z� /       malorum     l��fU  �l��fU  `m�sed do eiusmo tempo incidunt ut labore et dolor magna aliq    ����  ��� /       bonorum     p%��fU  0&��fU  �&�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  "����  ��� /       bonorum tion B��fU  PY��fU  �D�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  #����  ��� /       bonorum tion E��fU  pF��fU  0G�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  $����  ��� /       bonorum tion ��fU  ���fU  0�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �{���  ��� /      bonorum     �X��fU  pY��fU  0Z�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��"��  CŴ /       exercitation                   Lorem ipsum dolor sit amet, consectetur adipiscing elit      ��"��  CŴ /       exercitation ���fU  й��fU  P��Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  ��"��  CŴ /       exercitation ���fU   ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  ��"��  CŴ /       exercitation ���fU  ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  p],��  �Ǵ /       Birthday                       ullamco laboris nisi ut aliquip ex ea commodo consequat      s],��  �Ǵ /       Birthday    P��fU  ��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  u],��  �Ǵ /       Birthday     ��fU  ���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  w],��  �Ǵ /       Birthday    @*��fU  �*��fU  �+�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  v:��  J˴ /      exercitation                   Duis aute irure dolor in rehendert in volupate velit esse    `����  �� /       consectetur ����fU  @���fU  ���cillum dolore eu fugiat nulla pariatur  adipiscing elit �fU  a����  �� /       consectetur �I��fU  @J��fU  �J�cillum dolore eu fugiat nulla pariatur  adipiscing elit �fU  ��^��  8� /       Workout     B��fU  pL��fU  �C�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��^��  8� /       Workout fU  ����fU  ����fU  @��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��^��  8� /       Workout     ����fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��^��  8� /       Workout     ����fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �C���  0e� /       Workout fU  ����fU  �	��fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  �C���  0e� /       Workout     0���fU  ����fU  0��sunt in culpa qui offici desunt molit aim id est laborum. U  �C���  0e� /       Workout     0���fU  ����fU  0��sunt in culpa qui offici desunt molit aim id est laborum. U  �C���  0e� /       Workout fU  P\��fU  �\��fU  P]�sunt in culpa qui offici desunt molit aim id est laborum. U  d:��  @�� /      Appointment ����fU  ����fU  p��Duis aute irure dolor in rehendert in volupate velit esse U  I����  }�� /       Appointment @���fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  J����  }�� /       Appointment  ���fU  `���fU   ��Duis aute irure dolor in rehendert in volupate velit esse    �����  1�� /      exercitation 6��fU  �6��fU  �7�Duis aute irure dolor in rehendert in volupate velit esse U  �#F��  �Ե /       Appointment `j��fU  �j��fU  �v�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �#F��  �Ե /       Appointment �i��fU  j��fU  �j�ullamco laboris nisi ut aliquip ex ea commodo consequat iq   �#F��  �Ե /       Appointment ����fU  ���fU  Ч�ullamco laboris nisi ut aliquip ex ea commodo consequat iq   �#F��  �Ե /       Appointment �\��fU  �^��fU  b�ullamco laboris nisi ut aliquip ex ea commodo consequat iq   m�b��  �۵ /      bonorum     0T��fU  �T��fU  pU�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  @Zx��  �"� /       Birthday    ����fU   ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  AZx��  �"� /       Birthday    `r��fU  s��fU  �s�Duis aute irure dolor in rehendert in volupate velit esse U   ?���  �p� /       exercitation @��fU  A��fU  �A�Duis aute irure dolor in rehendert in volupate velit esse U  !?���  �p� /       exercitation Q��fU  �Q��fU   R�Duis aute irure dolor in rehendert in volupate velit esse U  "?���  �p� /       exercitation L��fU  @M��fU   N�Duis aute irure dolor in rehendert in volupate velit esse U  #?���  �p� /       exercitation 9��fU  @C��fU  �:�Duis aute irure dolor in rehendert in volupate velit esse U  ��A��  �� /       Birthday ur ���fU  ���fU  �ullamco laboris nisi ut aliquip ex ea commodo consequat e U  ��A��  �� /       Birthday ur  ��fU   ��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat e U  HG��  ]�� /       bonorum fU  `���fU   ���fU  ���cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  JG��  ]�� /       bonorum     �"��fU  p#��fU  �#�cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  KG��  ]�� /       bonorum     ���fU   ��fU  ��cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  MG��  ]�� /       bonorum     ���fU  @��fU   �cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  ]+a��  �� /      Birthday    <��fU  �<��fU  �=�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ^���  ��� /       consectetur                    sed do eiusmo tempo incidunt ut labore et dolor magna aliq   
^���  ��� /       consectetur �@��fU  PA��fU  B�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ^���  ��� /       consectetur P���fU  й��fU  P��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ^���  ��� /       consectetur 0���fU  ����fU  0��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �����  �¶ /       Birthday    �]��fU  0^��fU  �^�Duis aute irure dolor in rehendert in volupate velit esse U  �����  �¶ /       Birthday    p���fU  ����fU  � �Duis aute irure dolor in rehendert in volupate velit esse U  1����  ^ƶ /       Birthday U  ����fU  `���fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  3����  ^ƶ /       Birthday    0v��fU  �v��fU  pw�Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   5����  ^ƶ /       Birthday    �u��fU  0v��fU  �v�Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   8����  ^ƶ /       Birthday U  PE��fU  �E��fU  �F�Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   ��iq,�  �\ &/      malorum fU  ����fU  ����fU  @��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��tq,�  d_ &/       malorum                        cillum dolore eu fugiat nulla pariatur                       ��tq,�  d_ &/       malorum     ���fU  P��fU  �cillum dolore eu fugiat nulla pariatur ��fU  0��fU  ���fU  ��tq,�  d_ &/       malorum     �z��fU  �{��fU  p|�cillum dolore eu fugiat nulla pariatur ��fU  ����fU  p���fU  ��tq,�  d_ &/       malorum     P\��fU  �\��fU  �]�cillum dolore eu fugiat nulla pariatur ��fU  �`��fU  0a��fU  -vq,�  �_ &/       exercitation ^��fU  �^��fU  _�Excepteur sint occaecat cupidatat non proident ��fU  �c��fU  -vq,�  �_ &/       exercitation ���fU  ����fU  @��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �׀q,�  �b &/       exercitation ��fU   ��fU  ��Excepteur sint occaecat cupidatat non proident ��fU  �!��fU  �׀q,�  �b &/       exercitation ���fU  ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  P���fU  �׀q,�  �b &/       exercitation ��fU  ��fU  ��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  �׀q,�  �b &/       exercitation ���fU  0���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  `���fU  ��r,�  � &/      Birthday U  `��fU  ���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  Tsut,�  6$&/      bonorum     p���fU  0���fU  ���Excepteur sint occaecat cupidatat non proident onsequat �fU  �M�u,�  �n&/       exercitation x��fU  py��fU  0}�Excepteur sint occaecat cupidatat non proident ��fU  Ћ��fU  �M�u,�  �n&/       exercitation ���fU  ����fU   ��Excepteur sint occaecat cupidatat non proident ��fU   ���fU  �M�u,�  �n&/       exercitation ���fU  ����fU  P��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �M�u,�  �n&/       exercitation C��fU  @D��fU  00�Excepteur sint occaecat cupidatat non proident ��fU  �4��fU  ;��u,�  Sr&/       malorum     ���fU  ����fU  ��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  =��u,�  Sr&/       malorum     �h��fU  @i��fU  �i�Excepteur sint occaecat cupidatat non proident ��fU  ���fU  �=6v,�  �&/       Workout     �x��fU  py��fU  0}�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �=6v,�  �&/       Workout     ���fU  `���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �=6v,�  �&/       Workout     ����fU  @���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �=6v,�  �&/       Workout fU  ����fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU   <v,�  ��&/       Birthday                       Lorem ipsum dolor sit amet, consectetur adipiscing elit      #<v,�  ��&/       Birthday    P7��fU  �7��fU  �8�Lorem ipsum dolor sit amet, consectetur adipiscing elit e    &<v,�  ��&/       Birthday    `s��fU   t��fU  �t�Lorem ipsum dolor sit amet, consectetur adipiscing elit e    )<v,�  ��&/       Birthday U  ����fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit e    2�=v,�  ��&/       malorum tur ����fU  ����fU  @��cillum dolore eu fugiat nulla pariatur ommodo consequat . U  5�=v,�  ��&/       malorum tur `r��fU   s��fU  �s�cillum dolore eu fugiat nulla pariatur ommodo consequat .    8�=v,�  ��&/       malorum tur �C��fU  @D��fU   E�cillum dolore eu fugiat nulla pariatur ommodo consequat .    ;�=v,�  ��&/       malorum tur �t��fU  u��fU   v�cillum dolore eu fugiat nulla pariatur ommodo consequat .    ��v,�  +�&/       Birthday    p���fU  ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  ��v,�  +�&/       Birthday     ���fU  ����fU   ��sunt in culpa qui offici desunt molit aim id est laborum. U  <l�v,�  W�&/      malorum fU  p���fU  0���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �Mdw,�  n�&/       bonorum fU  �M��fU   N��fU   Q�Duis aute irure dolor in rehendert in volupate velit esse U  �Mdw,�  n�&/       bonorum ent ����fU  0���fU  ���Duis aute irure dolor in rehendert in volupate velit esse    �Mdw,�  n�&/       bonorum ent ����fU  ����fU   ��Duis aute irure dolor in rehendert in volupate velit esse    �Mdw,�  n�&/       bonorum ent ����fU  p���fU  0��Duis aute irure dolor in rehendert in volupate velit esse    |��w,�  _
&/      bonorum fU  ���fU  P��fU  �Excepteur sint occaecat cupidatat non proident ��fU  ���fU  q��w,�  f&/       Workout     �+��fU  ,��fU  �,�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  r��w,�  f&/       Workout     0���fU  ����fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  䲍x,�  �0&/      malorum                        Duis aute irure dolor in rehendert in volupate velit esse    �y8y,�  H\&/      bonorum                        Duis aute irure dolor in rehendert in volupate velit esse    X½y,�  g~&/       Birthday                       sunt in culpa qui offici desunt molit aim id est laborum.    Z½y,�  g~&/       Birthday    � ��fU  P!��fU  �!�sunt in culpa qui offici desunt molit aim id est laborum. U  [½y,�  g~&/       Birthday    p(��fU  0)��fU  0*�sunt in culpa qui offici desunt molit aim id est laborum. U  \½y,�  g~&/       Birthday    �8��fU  `9��fU   :�sunt in culpa qui offici desunt molit aim id est laborum. U  UU�y,�  v�&/      Meeting     �7��fU  `8��fU   9�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ���z,�  3�&/      Birthday    ����fU  `���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  H��{,�  }�&/       Workout     �C��fU  @D��fU   E�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  I��{,�  }�&/       Workout     0&��fU  �&��fU  0'�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  <�0|,�  �&/      bonorum                        Duis aute irure dolor in rehendert in volupate velit esse    ��|,�  �F&/      bonorum fU  ����fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �*�|,�  6G&/       malorum     p^��fU  0_��fU  �_�Duis aute irure dolor in rehendert in volupate velit esse U  �*�|,�  6G&/       malorum     `���fU  ����fU  `��Duis aute irure dolor in rehendert in volupate velit esse U  �*�|,�  6G&/       malorum     ����fU  ����fU  `��Duis aute irure dolor in rehendert in volupate velit esse U  �*�|,�  6G&/       malorum     �&��fU  p'��fU  �)�Duis aute irure dolor in rehendert in volupate velit esse U  �R},�  �h&/      Meeting     �&��fU  p'��fU  �)�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ���,�  �&/      consectetur P@��fU  A��fU  �A�Duis aute irure dolor in rehendert in volupate velit esse U  �ּ,�  b&/       bonorum     ����fU  P���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �ּ,�  b&/       bonorum ent                    ullamco laboris nisi ut aliquip ex ea commodo consequat e    �ּ,�  b&/       bonorum ent �b��fU  c��fU  �c�ullamco laboris nisi ut aliquip ex ea commodo consequat e U  �ּ,�  b&/       bonorum ent  ��fU  ���fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat e U  `0�,�  �&/       Appointment ����fU  ����fU  @��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  ����fU  c0�,�  �&/       Appointment  H��fU   I��fU  �I�cillum dolore eu fugiat nulla pariatur ommodo consequat e U  e0�,�  �&/       Appointment  4��fU   5��fU  �5�cillum dolore eu fugiat nulla pariatur ommodo consequat e U  g0�,�  �&/       Appointment  t��fU   u��fU  �u�cillum dolore eu fugiat nulla pariatur ommodo consequat e U  ��Y�,�  �/&/      Meeting fU  P
��fU  �
��fU  ��cillum dolore eu fugiat nulla pariatur ��fU  ���fU  ��fU  мg�,�  "3&/       Birthday    @���fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  Ҽg�,�  "3&/       Birthday ion ��fU  ���fU  P�ullamco laboris nisi ut aliquip ex ea commodo consequat . U  Ӽg�,�  "3&/       Birthday ion V��fU  �V��fU  �L�ullamco laboris nisi ut aliquip ex ea commodo consequat . U  Լg�,�  "3&/       Birthday ion ��fU  ��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat . U  �G��,�  ^W&/      Appointment                    sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��$�,�  �&/      bonorum     0���fU  ���fU  p��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ���,�  .�&/       Appointment P6��fU  �6��fU  P7�Duis aute irure dolor in rehendert in volupate velit esse U  ���,�  .�&/       Appointment ����fU   ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse    ���,�  .�&/       Appointment ����fU  @���fU  ���Duis aute irure dolor in rehendert in volupate velit esse    ���,�  .�&/       Appointment  ���fU  ����fU   ��Duis aute irure dolor in rehendert in volupate velit esse    4��,�  �&/      Birthday    P��fU  ��fU  `�sunt in culpa qui offici desunt molit aim id est laborum. U  쨱�,�  !�&/       consectetur ���fU  �	��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �,�  !�&/       consectetur P���fU  ����fU  P��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��g�,�  �v&/      Meeting     p��fU  0��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  ��~�,�  �|&/       malorum     ����fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ±~�,�  �|&/       malorum     �}��fU   ~��fU  �~�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �g�,�  V�&/       bonorum     p���fU  0���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  `���fU  �g�,�  V�&/       bonorum     p���fU  0���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  P���fU  �g�,�  V�&/       bonorum      ���fU  ����fU  0��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �g�,�  V�&/       bonorum     '��fU  �'��fU  P(�Excepteur sint occaecat cupidatat non proident ��fU  -��fU  K��,�  ��&/      Appointment pw��fU  �w��fU  px�sunt in culpa qui offici desunt molit aim id est laborum. U  ,AѮ,�  �&/      Birthday     	��fU  ��fU  P
�sunt in culpa qui offici desunt molit aim id est laborum. U  �e�,�  �:&/       Workout     �>��fU   ?��fU  �?�Excepteur sint occaecat cupidatat non proident ��fU  `C��fU  �e�,�  �:&/       Workout     ���fU  ����fU  0��Excepteur sint occaecat cupidatat non proident ��fU  О��fU  99h�,�  s;&/       Birthday    ����fU  @���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ;9h�,�  s;&/       Birthday    `���fU  ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   D m�,�  �<&/      Workout                        Excepteur sint occaecat cupidatat non proident               <e
�,�  �d&/      Meeting     �&��fU  p'��fU  �)�Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  1z�,�  >e&/       malorum     P,��fU  -��fU  �-�cillum dolore eu fugiat nulla pariatur ��fU  P1��fU  �1��fU  2z�,�  >e&/       malorum     �{��fU   |��fU  �|�cillum dolore eu fugiat nulla pariatur ��fU   ���fU  ����fU  �`$�,�  '�&/      Meeting                        sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �o5�,�  ��&/       Birthday U  0���fU   ���fU  P��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �o5�,�  ��&/       Birthday    ����fU   ���fU  P��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �o5�,�  ��&/       Birthday    ����fU  ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �o5�,�  ��&/       Birthday    p���fU  ����fU  p��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �T��,�  O�&/       Workout      ���fU  ����fU  0��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �T��,�  O�&/       Workout     ����fU  `���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��,�  �(&/      Birthday    �[��fU  0\��fU  �\�cillum dolore eu fugiat nulla pariatur ��fU  `��fU  �`��fU  �r�,�  a+&/       exercitation X��fU  pY��fU  0Z�sunt in culpa qui offici desunt molit aim id est laborum. U  �r�,�  a+&/       exercitation 	��fU  p
��fU   �sunt in culpa qui offici desunt molit aim id est laborum.    �r�,�  a+&/       exercitation )��fU  *��fU  �*�sunt in culpa qui offici desunt molit aim id est laborum.    �r�,�  a+&/       exercitation ���fU  `���fU  ���sunt in culpa qui offici desunt molit aim id est laborum.    Xї�,�  �M&/       Workout tion 5��fU  `6��fU  �6�Excepteur sint occaecat cupidatat non proident  magna aliq   Yї�,�  �M&/       Workout tion 4��fU  �4��fU  P5�Excepteur sint occaecat cupidatat non proident  magna aliq   4Է�,�  ��&/      Appointment @���fU   ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  yXǴ,�  {�&/       Birthday ion ���fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  zXǴ,�  {�&/       Birthday ion w��fU  `x��fU  �x�Duis aute irure dolor in rehendert in volupate velit esse    {XǴ,�  {�&/       Birthday ion x��fU  0y��fU  �y�Duis aute irure dolor in rehendert in volupate velit esse    |XǴ,�  {�&/       Birthday ion t��fU  �u��fU   ��Duis aute irure dolor in rehendert in volupate velit esse    d�h�,�  ��&/      malorum tur ����fU  ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   �	�,�  ��&/       Appointment                    cillum dolore eu fugiat nulla pariatur                       �	�,�  ��&/       Appointment  c��fU  �c��fU  �d�cillum dolore eu fugiat nulla pariatur et dolor magna aliq   �	�,�  ��&/       Appointment ����fU   ���fU  ���cillum dolore eu fugiat nulla pariatur et dolor magna aliq   �	�,�  ��&/       Appointment @���fU   ���fU  ���cillum dolore eu fugiat nulla pariatur et dolor magna aliq   ���,�  e�&/       malorum ent ����fU  ����fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  ���,�  e�&/       malorum ent ���fU  p��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  ���,�  e�&/       malorum ent ����fU  ����fU  P��Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  ���,�  e�&/       malorum ent P��fU  ���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  ���,�  &/      consectetur                    sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ԓ��,�  �&/       consectetur  f��fU  �f��fU  �g�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ֓��,�  �&/       consectetur  J��fU  �J��fU   K�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  iE��,�  �&/       Workout fU  0���fU  ����fU  p��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   jE��,�  �&/       Workout ent ����fU  ����fU  @��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   kE��,�  �&/       Workout ent ����fU  @���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   mE��,�  �&/       Workout ent  ���fU  ����fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   4~Z�,�  &/      exercitation &��fU  p'��fU  �)�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   QDn�,�  Ҋ&/       malorum     P���fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  RDn�,�  Ҋ&/       malorum fU  `��fU  ���fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �惹,�  ��&/      exercitation ���fU  ����fU  `��sunt in culpa qui offici desunt molit aim id est laborum. U   &��,�  �&/       malorum fU  U��fU  �U��fU  Y�cillum dolore eu fugiat nulla pariatur ��fU  @f��fU   g��fU  !&��,�  �&/       malorum tion [��fU  0\��fU  �\�cillum dolore eu fugiat nulla pariatur et dolor magna aliq   "&��,�  �&/       malorum tion ���fU   ���fU  ���cillum dolore eu fugiat nulla pariatur et dolor magna aliq   $&��,�  �&/       malorum tion ���fU  ����fU   ��cillum dolore eu fugiat nulla pariatur et dolor magna aliq   �!�,�  Y�&/      malorum fU  ����fU  ����fU  @��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   h;˺,�  �%&/       Meeting fU  p���fU  0���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  i;˺,�  �%&/       Meeting fU  ����fU  ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  j;˺,�  �%&/       Meeting     �8��fU  �9��fU  :�sunt in culpa qui offici desunt molit aim id est laborum. U  k;˺,�  �%&/       Meeting     `<��fU   =��fU  �=�sunt in culpa qui offici desunt molit aim id est laborum. U  Х�,�  �n&/       Appointment �1��fU  �2��fU  `3�Excepteur sint occaecat cupidatat non proident ��fU  `8��fU  ѥ�,�  �n&/       Appointment 0���fU  ���fU  p��Excepteur sint occaecat cupidatat non proident onsequat �fU  ҥ�,�  �n&/       Appointment D��fU  �D��fU  �G�Excepteur sint occaecat cupidatat non proident onsequat �fU  ӥ�,�  �n&/       Appointment `���fU  ���fU  `��Excepteur sint occaecat cupidatat non proident onsequat �fU  ���,�  g�&/      bonorum     0���fU  ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ���,�  d�&/      Meeting     ����fU  P ��fU  � �sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ���,�  �/&/      Meeting     p��fU  0��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��b�,�  �T&/       consectetur  ���fU  ����fU  `��sunt in culpa qui offici desunt molit aim id est laborum. U  ��b�,�  �T&/       consectetur ����fU  p���fU  0��sunt in culpa qui offici desunt molit aim id est laborum. U  ��b�,�  �T&/       consectetur px��fU  0y��fU  �y�sunt in culpa qui offici desunt molit aim id est laborum. U  ��b�,�  �T&/       consectetur Ѝ��fU  P���fU   ��sunt in culpa qui offici desunt molit aim id est laborum. U  #Vd�,�  U&/       Appointment �7��fU  `8��fU   9�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  %Vd�,�  U&/       Appointment `���fU  ���fU  `��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��,�  ��&/      bonorum     D��fU  �D��fU  �G�Duis aute irure dolor in rehendert in volupate velit esse U  ��,�  ?�&/       Meeting fU  ����fU  ����fU  @��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  `���fU  ��,�  ?�&/       Meeting     ���fU  p���fU  ��cillum dolore eu fugiat nulla pariatur ��fU  @���fU  ����fU  o9��,�  u�&/      bonorum     ����fU   ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  躩�,�  a�&/       exercitation ��fU  ���fU  � �sunt in culpa qui offici desunt molit aim id est laborum. U  麩�,�  a�&/       exercitation &��fU  p'��fU  �)�sunt in culpa qui offici desunt molit aim id est laborum. U  꺩�,�  a�&/       exercitation ���fU  ����fU  @��sunt in culpa qui offici desunt molit aim id est laborum. U  캩�,�  a�&/       exercitation ���fU  ����fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  $���,�  ��&/      exercitation ���fU   ���fU  P��ullamco laboris nisi ut aliquip ex ea commodo consequat e U  ���,�  ��&/       Appointment P��fU  ��fU  0/�cillum dolore eu fugiat nulla pariatur ��fU  P��fU  ���fU  ���,�  ��&/       Appointment ����fU  `���fU   ��cillum dolore eu fugiat nulla pariatur ��fU  `���fU   ���fU  ���,�  ��&/       Appointment ����fU  ����fU  `��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  ����fU  ���,�  ��&/       Appointment ����fU  P���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ���fU  P��fU  �,b�,�  " &/       Workout     �9��fU  P:��fU  �1�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �,b�,�  " &/       Workout     D��fU  �D��fU  �G�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �,b�,�  " &/       Workout     ����fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �,b�,�  " &/       Workout     @���fU  ����fU  @��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��,�  �C &/      Meeting     <��fU  �<��fU  �=�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ���,�  j &/       Birthday    ��fU  ���fU  P�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ���,�  j &/       Birthday    ���fU  0 ��fU  � �Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �&�,�  Ќ &/       bonorum     ���fU  ���fU  p�cillum dolore eu fugiat nulla pariatur ��fU  @��fU   ��fU  �&�,�  Ќ &/       bonorum     ����fU  ����fU  P��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  ����fU  �&�,�  Ќ &/       bonorum     p���fU  ����fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU  P���fU  �&�,�  Ќ &/       bonorum     ?��fU  �?��fU  P@�cillum dolore eu fugiat nulla pariatur ��fU  �D��fU  @E��fU  }F;�,�  ?� &/      consectetur P���fU  ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   !h��,�  T� &/       exercitation ���fU  ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  "h��,�  T� &/       exercitation X��fU  �X��fU  `Y�sunt in culpa qui offici desunt molit aim id est laborum. U  D���,�  ̻ &/      Birthday    U��fU  �U��fU  Y�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��p�,�  �� &/       malorum     ����fU  ����fU  @��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  ��p�,�  �� &/       malorum     b��fU  �b��fU  Pc�Excepteur sint occaecat cupidatat non proident ��fU  �g��fU  ��p�,�  �� &/       malorum                        Excepteur sint occaecat cupidatat non proident               ��p�,�  �� &/       malorum     ����fU  P���fU  Ќ�Excepteur sint occaecat cupidatat non proident ��fU  ����fU  ,�s�,�  M� &/      Appointment ����fU  P���fU  ��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  ���,�  a!&/       Workout                        Lorem ipsum dolor sit amet, consectetur adipiscing elit      ���,�  a!&/       Workout     ��fU  ���fU  P�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ���,�  a!&/       Workout     �w��fU  `x��fU  �x�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ���,�  a!&/       Workout     ���fU  ���fU  p�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ����,�  !&/      Workout                        Lorem ipsum dolor sit amet, consectetur adipiscing elit      Z��,�  '!&/       Appointment  ��fU  ���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  \��,�  '!&/       Appointment ����fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ^��,�  '!&/       Appointment                    Lorem ipsum dolor sit amet, consectetur adipiscing elit      `��,�  '!&/       Appointment 0���fU  ����fU  p��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  x[��,�  [+!&/       Birthday    ���fU  ����fU  ��cillum dolore eu fugiat nulla pariatur ��fU  @���fU  ����fU  y[��,�  [+!&/       Birthday    ����fU   ���fU  ���cillum dolore eu fugiat nulla pariatur ��fU   ��fU  ���fU  �x��,�  )w!&/      Birthday U  ����fU  ����fU  @��Excepteur sint occaecat cupidatat non proident ��fU  `���fU  4�M�,�  "�!&/      Appointment                    Duis aute irure dolor in rehendert in volupate velit esse    Dc��,�  ��!&/      Birthday                       Duis aute irure dolor in rehendert in volupate velit esse    ���,�  7�!&/       consectetur D��fU  �D��fU  �G�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ���,�  7�!&/       consectetur ����fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ���,�  �"&/       Birthday     ���fU  ����fU   x�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ���,�  �"&/       Birthday    0.��fU  �.��fU  `/�ullamco laboris nisi ut aliquip ex ea commodo consequat e U  ����,�  (?"&/      exercitation D��fU  �D��fU  �G�cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  �Gj�,�  i"&/      bonorum     �&��fU  p'��fU  �)�Excepteur sint occaecat cupidatat non proident ��fU  �5��fU  W��,�  �"&/      Birthday    p���fU  0���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  � �,�  ��"&/       bonorum                        Duis aute irure dolor in rehendert in volupate velit esse    
� �,�  ��"&/       bonorum     ���fU  и��fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  � �,�  ��"&/       bonorum     ���fU  ���fU   �Duis aute irure dolor in rehendert in volupate velit esse U  � �,�  ��"&/       bonorum     ����fU  ����fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  �� �,�  9�"&/       bonorum                        Excepteur sint occaecat cupidatat non proident               �� �,�  9�"&/       bonorum     V��fU  �V��fU  �L�Excepteur sint occaecat cupidatat non proident ��fU  �Q��fU  �� �,�  9�"&/       bonorum     ����fU  P���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ���fU  �� �,�  9�"&/       bonorum fU  0���fU  Н��fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  y�$�,�  [�"&/       Birthday    �x��fU  py��fU  0}�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   {�$�,�  [�"&/       Birthday    @f��fU   g��fU  �j�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   }�$�,�  [�"&/       Birthday    ����fU  `���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �$�,�  [�"&/       Birthday    p���fU  ���fU  p��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �|W�,�  �(#&/      Workout                        Duis aute irure dolor in rehendert in volupate velit esse    Q�e�,�  r,#&/       Appointment ����fU  P���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  R�e�,�  r,#&/       Appointment `��fU  ���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  S�e�,�  r,#&/       Appointment ����fU   ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  T�e�,�  r,#&/       Appointment �A��fU  @B��fU  �B�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ���,�  �S#&/      exercitation ���fU  `���fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  `p�$-�  �O.&/       Appointment 0���fU  ����fU  p��Excepteur sint occaecat cupidatat non proident ��fU  0���fU  ap�$-�  �O.&/       Appointment 0	��fU  �	��fU  0
�Excepteur sint occaecat cupidatat non proident ��fU   ��fU  bp�$-�  �O.&/       Appointment ����fU  `���fU   ��Excepteur sint occaecat cupidatat non proident ��fU  `���fU  cp�$-�  �O.&/       Appointment p���fU  0���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  0���fU  �^%-�  Nn.&/      Meeting     0J��fU  �J��fU  0K�sunt in culpa qui offici desunt molit aim id est laborum. U  �l%-�  �q.&/       consectetur `���fU  ���fU  `��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  �l%-�  �q.&/       consectetur ����fU  `���fU  ���Excepteur sint occaecat cupidatat non proident onsequat .    �&�%-�  ��.&/       Birthday U  0���fU  ����fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  �&�%-�  ��.&/       Birthday    _��fU  �_��fU  �`�sunt in culpa qui offici desunt molit aim id est laborum. U  �&�%-�  ��.&/       Birthday    p(��fU  0)��fU  0*�sunt in culpa qui offici desunt molit aim id est laborum. U  �&�%-�  ��.&/       Birthday    a��fU  �a��fU  pb�sunt in culpa qui offici desunt molit aim id est laborum. U  J&-�  ��.&/       Workout     ����fU  @���fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  J&-�  ��.&/       Workout      c��fU  �c��fU   d�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  |2&-�  ��.&/      Workout fU  �x��fU  py��fU  0}�sunt in culpa qui offici desunt molit aim id est laborum. U  ��&-�  �.&/      Birthday    ���fU  P���fU  Ѐ�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ���&-�  y�.&/       exercitation _��fU  @`��fU  �`�Excepteur sint occaecat cupidatat non proident ��fU  �d��fU  ���&-�  y�.&/       exercitation ��fU  ���fU  ��Excepteur sint occaecat cupidatat non proident ��fU   ��fU  �&-�  U�.&/       malorum     ��fU  ���fU  P�cillum dolore eu fugiat nulla pariatur ��fU  ��fU  ���fU  �&-�  U�.&/       malorum      '��fU  �'��fU  P(�cillum dolore eu fugiat nulla pariatur ��fU  �+��fU  PM��fU  9�.'-�  �.&/       Appointment                    sed do eiusmo tempo incidunt ut labore et dolor magna aliq   :�.'-�  �.&/       Appointment ���fU  Ћ��fU  Џ�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ;�.'-�  �.&/       Appointment P5��fU  �5��fU  P6�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   <�.'-�  �.&/       Appointment 0)��fU  �)��fU  0*�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   \e;'-�  K�.&/      consectetur                    Duis aute irure dolor in rehendert in volupate velit esse    �'-�  �/&/      malorum     �!��fU  P"��fU  #�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  $i�)-�  ��/&/      bonorum fU  ���fU  P��fU  �sunt in culpa qui offici desunt molit aim id est laborum. U  9�)-�  ��/&/       exercitation <��fU  �<��fU  �=�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  :�)-�  ��/&/       exercitation ��fU  ���fU  p�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ;�)-�  ��/&/       exercitation ��fU  @��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  <�)-�  ��/&/       exercitation _��fU  �_��fU  �`�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �zB*-�  ��/&/       exercitation ��fU   ��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  �zB*-�  ��/&/       exercitation ���fU  ���fU  `��sunt in culpa qui offici desunt molit aim id est laborum. U  X��*-�  ��/&/       Appointment P���fU  ���fU  У�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  Z��*-�  ��/&/       Appointment ����fU   ���fU  P��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  [��*-�  ��/&/       Appointment  ���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  \��*-�  ��/&/       Appointment @���fU  ����fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��*-�  ��/&/      Meeting     �t��fU  �u��fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �?\+-�  ��/&/       Appointment                    Duis aute irure dolor in rehendert in volupate velit esse    �?\+-�  ��/&/       Appointment P
��fU  �
��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  �?\+-�  ��/&/       Appointment �@��fU  PA��fU  B�Duis aute irure dolor in rehendert in volupate velit esse U  �?\+-�  ��/&/       Appointment ����fU    ��fU  � �Duis aute irure dolor in rehendert in volupate velit esse U  <0,-�  �!0&/      exercitation R��fU  pS��fU  0T�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �V�,-�  �F0&/      Meeting     ����fU   ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  X}�--�  G�0&/       Meeting     �t��fU  �u��fU   ��sunt in culpa qui offici desunt molit aim id est laborum. U  [}�--�  G�0&/       Meeting     @���fU  ����fU  @��sunt in culpa qui offici desunt molit aim id est laborum. U  ]}�--�  G�0&/       Meeting     ����fU  P���fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  _}�--�  G�0&/       Meeting     �n��fU   o��fU  �o�sunt in culpa qui offici desunt molit aim id est laborum. U  ��--�  ��0&/      Birthday    ���fU  ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  2��--�  >�0&/       consectetur P���fU  ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  4��--�  >�0&/       consectetur ����fU  ����fU  P��sunt in culpa qui offici desunt molit aim id est laborum. U  6��--�  >�0&/       consectetur p���fU   ���fU   ��sunt in culpa qui offici desunt molit aim id est laborum. U  8��--�  >�0&/       consectetur  ��fU  ���fU   �sunt in culpa qui offici desunt molit aim id est laborum. U  ̊b.-�  �0&/      malorum     ����fU   ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �M/-�  E�0&/       bonorum     ���fU  н��fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU  P���fU  �M/-�  E�0&/       bonorum  ion O��fU  �P��fU   Q�cillum dolore eu fugiat nulla pariatur roident ing elit e    �M/-�  E�0&/       bonorum  ion M��fU  PN��fU  �N�cillum dolore eu fugiat nulla pariatur roident ing elit e    �M/-�  E�0&/       bonorum  ion V��fU  �V��fU  0W�cillum dolore eu fugiat nulla pariatur roident ing elit e     ڗ/-�  @1&/       Appointment `��fU  �`��fU  Pa�sunt in culpa qui offici desunt molit aim id est laborum. U  ڗ/-�  @1&/       Appointment  ���fU  ����fU  @��sunt in culpa qui offici desunt molit aim id est laborum. U  � �0-�  �V1&/      Workout     @���fU   ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ��P1-�  }1&/       exercitation r��fU  Ps��fU  �s�Excepteur sint occaecat cupidatat non proident ��fU  Pw��fU  ��P1-�  }1&/       exercitation ���fU  @���fU  ���Excepteur sint occaecat cupidatat non proident onsequat �fU  <�a1-�  w�1&/      bonorum                        Excepteur sint occaecat cupidatat non proident               -�1-�  $�1&/      exercitation                   ullamco laboris nisi ut aliquip ex ea commodo consequat      �E�1-�  �1&/       Birthday nt �9��fU  P:��fU  �1�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �E�1-�  �1&/       Birthday nt ����fU  ���fU  л�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �E�1-�  �1&/       Birthday nt                    ullamco laboris nisi ut aliquip ex ea commodo consequat      �E�1-�  �1&/       Birthday nt p���fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �2-�  ?�1&/      Meeting      ��fU  ���fU  P�Duis aute irure dolor in rehendert in volupate velit esse U  &�2-�  ��1&/       consectetur @���fU   ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  	&�2-�  ��1&/       consectetur 0���fU  ����fU  p��Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  
&�2-�  ��1&/       consectetur                    Lorem ipsum dolor sit amet, consectetur adipiscing elit .    &�2-�  ��1&/       consectetur P���fU  ����fU  P��Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  8d3-�  ��1&/      consectetur ����fU  ����fU  @��sunt in culpa qui offici desunt molit aim id est laborum. U  �,3-�  ��1&/       malorum fU   H��fU  �H��fU  �I�Duis aute irure dolor in rehendert in volupate velit esse U  �,3-�  ��1&/       malorum     ����fU  ����fU  `��Duis aute irure dolor in rehendert in volupate velit esse U  �,3-�  ��1&/       malorum     �+��fU  p,��fU  �,�Duis aute irure dolor in rehendert in volupate velit esse U  �,3-�  ��1&/       malorum fU  g��fU  ����fU  =�Duis aute irure dolor in rehendert in volupate velit esse U  PT$3-�  ��1&/       Workout tion                   sed do eiusmo tempo incidunt ut labore et dolor magna aliq   UT$3-�  ��1&/       Workout tion ���fU   ���fU  P��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   YT$3-�  ��1&/       Workout tion D��fU  �D��fU  �G�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ^T$3-�  ��1&/       Workout tion ���fU  ����fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��)3-�  E�1&/       malorum fU  <��fU  �<��fU  �=�Duis aute irure dolor in rehendert in volupate velit esse U  ��)3-�  E�1&/       malorum     ����fU  `���fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  ��)3-�  E�1&/       malorum      ��fU  ���fU  � �Duis aute irure dolor in rehendert in volupate velit esse U  ��)3-�  E�1&/       malorum fU  ����fU  P���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  c303-�  ��1&/       malorum fU  0���fU  ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  h303-�  ��1&/       malorum fU  :��fU  �:��fU  ;�sunt in culpa qui offici desunt molit aim id est laborum. U  l303-�  ��1&/       malorum     ����fU  `���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  q303-�  ��1&/       malorum     �[��fU  0\��fU  �\�sunt in culpa qui offici desunt molit aim id est laborum. U  %�13-�  ?�1&/       Birthday    ����fU  p���fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  *�13-�  ?�1&/       Birthday    0���fU  ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �]�3-�  A2&/       Appointment                    sunt in culpa qui offici desunt molit aim id est laborum.    �]�3-�  A2&/       Appointment ?��fU  �?��fU  P@�sunt in culpa qui offici desunt molit aim id est laborum. U  �]�3-�  A2&/       Appointment �J��fU  �K��fU  V�sunt in culpa qui offici desunt molit aim id est laborum. U  �]�3-�  A2&/       Appointment `Y��fU  �Y��fU  �Z�sunt in culpa qui offici desunt molit aim id est laborum. U  ���3-�  �2&/      consectetur ����fU  `���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU   �H4-�  �?2&/       Appointment  ��fU  �!��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �H4-�  �?2&/       Appointment  d��fU  e��fU  �e�Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   �H4-�  �?2&/       Appointment  ���fU  @���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   �H4-�  �?2&/       Appointment  ���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   �]L4-�  �@2&/      Meeting      ��fU  ���fU  0�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �ZS4-�  eB2&/       Appointment ����fU   ���fU  ���cillum dolore eu fugiat nulla pariatur et dolor magna aliq   �ZS4-�  eB2&/       Appointment  ��fU  `��fU   �cillum dolore eu fugiat nulla pariatur et dolor magna aliq   5�g4-�  �G2&/       consectetur ����fU  0���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  8�g4-�  �G2&/       consectetur �5��fU  `6��fU  �6�Excepteur sint occaecat cupidatat non proident ��fU  �:��fU  p��4-�  &g2&/       exercitation ���fU  ����fU  P��Duis aute irure dolor in rehendert in volupate velit esse U  r��4-�  &g2&/       exercitation ���fU  ����fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  t��4-�  &g2&/       exercitation ���fU  @���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  v��4-�  &g2&/       exercitation ���fU  @���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ��4-�  *g2&/       Birthday nt ���fU  Ћ��fU  Џ�Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   ��4-�  *g2&/       Birthday nt ���fU  `��fU   	�Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   ��4-�  *g2&/       Birthday nt ����fU  ����fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   ��4-�  *g2&/       Birthday nt �"��fU  p#��fU  �#�Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   �K_-�  �B=&/      Appointment ���fU  P��fU  �cillum dolore eu fugiat nulla pariatur ��fU  0��fU  ���fU   w�_-�  �c=&/       Appointment @���fU  ����fU  @��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  !w�_-�  �c=&/       Appointment p���fU   ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  }��a-�  ?�=&/      exercitation ���fU  P ��fU  �ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��a-�  ��=&/       Workout fU  `���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  
��a-�  ��=&/       Workout     00��fU  �0��fU  P1�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��a-�  ��=&/       Workout fU  ���fU  0��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��a-�  ��=&/       Workout      c��fU  �c��fU   d�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �:b-�  �>&/       Workout     ����fU  `���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  	�:b-�  �>&/       Workout tur ����fU   ��fU   ��sunt in culpa qui offici desunt molit aim id est laborum. U  
�:b-�  �>&/       Workout tur � ��fU  �)��fU  p"�sunt in culpa qui offici desunt molit aim id est laborum. U  �:b-�  �>&/       Workout tur P��fU  ���fU  P�sunt in culpa qui offici desunt molit aim id est laborum. U  p d-�  �{>&/       malorum     ����fU  p���fU  P��Duis aute irure dolor in rehendert in volupate velit esse U  q d-�  �{>&/       malorum fU  0���fU  ����fU  0��Duis aute irure dolor in rehendert in volupate velit esse U  r d-�  �{>&/       malorum     0���fU  ����fU  p��Duis aute irure dolor in rehendert in volupate velit esse U  s d-�  �{>&/       malorum     p���fU  0���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  �Ѡd-�  ��>&/      bonorum fU  0��fU  ���fU  �	�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   $Ţd-�  t�>&/       malorum     p���fU  0���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  &Ţd-�  t�>&/       malorum      k��fU  �k��fU  Pl�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  	�d-�  �>&/       Birthday    �t��fU  �u��fU   ��sunt in culpa qui offici desunt molit aim id est laborum. U  
�d-�  �>&/       Birthday    �i��fU  j��fU  �j�sunt in culpa qui offici desunt molit aim id est laborum. U  �d-�  �>&/       Birthday    �e��fU  Pf��fU  g�sunt in culpa qui offici desunt molit aim id est laborum. U  �d-�  �>&/       Birthday    @|��fU  �|��fU  �}�sunt in culpa qui offici desunt molit aim id est laborum. U  ��e-�  ��>&/       consectetur P��fU  ��fU  `�Duis aute irure dolor in rehendert in volupate velit esse U  ��e-�  ��>&/       consectetur D��fU  �D��fU  �G�Duis aute irure dolor in rehendert in volupate velit esse U  ��e-�  ��>&/       consectetur ����fU  ����fU  `��Duis aute irure dolor in rehendert in volupate velit esse U  ��e-�  ��>&/       consectetur ����fU  0���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  3<`f-�  ~?&/       consectetur ���fU  �	��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  5<`f-�  ~?&/       consectetur  R��fU  �R��fU   S�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  H�df-�  �?&/       Appointment ����fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  I�df-�  �?&/       Appointment P���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  J�df-�  �?&/       Appointment ����fU  @���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  L�df-�  �?&/       Appointment @���fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  �!�f-�  �7?&/       Workout     ����fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �!�f-�  �7?&/       Workout     0���fU  ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  `-�f-�  8?&/       Birthday U  ����fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  b-�f-�  8?&/       Birthday    ����fU  P���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  c-�f-�  8?&/       Birthday    p���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  e-�f-�  8?&/       Birthday    @���fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��g-�  ??&/      bonorum     P���fU  ���fU  У�Excepteur sint occaecat cupidatat non proident ��fU  P���fU  ��g-�  �a?&/      Birthday    �&��fU  p'��fU  �)�cillum dolore eu fugiat nulla pariatur ��fU   5��fU  �5��fU  ��3h-�  +�?&/       consectetur �0��fU  `1��fU   5�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��3h-�  +�?&/       consectetur Ph��fU  �h��fU  �i�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��_i-�  ��?&/      Workout fU  `���fU  ����fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ,hj-�  -@&/      bonorum     ����fU  `���fU  ��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  ����fU  D9"k-�  LJ@&/      Birthday                       cillum dolore eu fugiat nulla pariatur                       �,�k-�  �o@&/      Workout                        sed do eiusmo tempo incidunt ut labore et dolor magna aliq   q�k-�  Fv@&/       Meeting     @f��fU   g��fU  �j�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  r�k-�  Fv@&/       Meeting     ����fU  0���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �pl-�  @&/       Meeting     ����fU  ����fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �pl-�  @&/       Meeting     `���fU   ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �pl-�  @&/       Meeting      ��fU  ���fU  0�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �pl-�  @&/       Meeting     ����fU  @���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  @C�l-�  ��@&/       Birthday U  0&��fU  �&��fU  0'�Excepteur sint occaecat cupidatat non proident ��fU  �*��fU  AC�l-�  ��@&/       Birthday    P)��fU  *��fU  �*�Excepteur sint occaecat cupidatat non proident ��fU  @D��fU  ��m-�  ��@&/      exercitation ���fU  ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  y%n-�  �A&/       bonorum     ����fU   ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  {%n-�  �A&/       bonorum ent �4��fU  `5��fU  �5�sunt in culpa qui offici desunt molit aim id est laborum. U  }%n-�  �A&/       bonorum ent P(��fU  �(��fU  P)�sunt in culpa qui offici desunt molit aim id est laborum. U  %n-�  �A&/       bonorum ent p��fU  0��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  01n-�  �A&/       bonorum     ����fU  p���fU  P��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  21n-�  �A&/       bonorum     � ��fU  P!��fU  �!�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  41n-�  �A&/       bonorum      '��fU  �'��fU  P(�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  61n-�  �A&/       bonorum     ���fU  ����fU  0��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  x�n-�  �5A&/       Workout                        Duis aute irure dolor in rehendert in volupate velit esse    y�n-�  �5A&/       Workout ent                    Duis aute irure dolor in rehendert in volupate velit esse    z�n-�  �5A&/       Workout ent `���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  {�n-�  �5A&/       Workout ent ����fU  `���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �
Ko-�  �ZA&/       Workout     ����fU  @���fU  P��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �
Ko-�  �ZA&/       Workout     0u��fU  �u��fU  0v�Excepteur sint occaecat cupidatat non proident ��fU  pz��fU  �
Ko-�  �ZA&/       Workout     ����fU  ����fU   ��Excepteur sint occaecat cupidatat non proident ��fU   ���fU  �
Ko-�  �ZA&/       Workout     ����fU  @���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �;�o-�  ځA&/       Appointment ����fU  p���fU  P��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �;�o-�  ځA&/       Appointment �#��fU  p$��fU  �$�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �;�o-�  ځA&/       Appointment px��fU  0y��fU  �y�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �;�o-�  ځA&/       Appointment ����fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ���o-�  Z�A&/       Appointment ��fU  ���fU  P�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ���o-�  Z�A&/       Appointment �r��fU  Ps��fU  �s�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  `*yp-�  <�A&/       Appointment                    sunt in culpa qui offici desunt molit aim id est laborum.    c*yp-�  <�A&/       Appointment  ���fU  @���fU   ��sunt in culpa qui offici desunt molit aim id est laborum. U  e*yp-�  <�A&/       Appointment  ��fU  @ ��fU  � �sunt in culpa qui offici desunt molit aim id est laborum. U  g*yp-�  <�A&/       Appointment  ��fU  �	��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  ��p-�  ��A&/      bonorum     P��fU  ��fU  `�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   )�p-�  �A&/       exercitation &��fU  p'��fU  �)�Excepteur sint occaecat cupidatat non proident ��fU  �5��fU  )�p-�  �A&/       exercitation ���fU  `���fU  ��Excepteur sint occaecat cupidatat non proident ��fU   ���fU  )�p-�  �A&/       exercitation ���fU  ����fU  @��Excepteur sint occaecat cupidatat non proident ��fU  `���fU   )�p-�  �A&/       exercitation ���fU  P���fU  ���Excepteur sint occaecat cupidatat non proident ��fU   ���fU  �q-�  ��A&/      Appointment ����fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �'�-�  /�L&/      bonorum     p���fU  0���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   D��-�  ��L&/      Appointment                    Lorem ipsum dolor sit amet, consectetur adipiscing elit      ���-�  ��L&/       consectetur D��fU  �D��fU  �G�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ���-�  ��L&/       consectetur @���fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  X�	�-�  G�L&/       Appointment                    Duis aute irure dolor in rehendert in volupate velit esse    Y�	�-�  G�L&/       Appointment ���fU  `��fU   	�Duis aute irure dolor in rehendert in volupate velit esse U  Z�	�-�  G�L&/       Appointment  ��fU  ���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  \�	�-�  G�L&/       Appointment � ��fU  `!��fU  "�Duis aute irure dolor in rehendert in volupate velit esse U  X/��-�  ��L&/       bonorum     p���fU  0���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  p���fU  Y/��-�  ��L&/       bonorum     �\��fU  �^��fU  b�Excepteur sint occaecat cupidatat non proident t laborum. U  Z/��-�  ��L&/       bonorum     ����fU  ���fU  ���Excepteur sint occaecat cupidatat non proident t laborum. U  [/��-�  ��L&/       bonorum     ����fU  @���fU  ���Excepteur sint occaecat cupidatat non proident t laborum. U  �J�-�  N!M&/       Workout                        sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �J�-�  N!M&/       Workout     0*��fU  �*��fU  �+�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �J�-�  N!M&/       Workout     `���fU   ���fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �J�-�  N!M&/       Workout     �u��fU  Pv��fU  �v�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��˝-�  �BM&/       malorum      ��fU  ���fU  � �cillum dolore eu fugiat nulla pariatur ��fU  p%��fU  0&��fU  ��˝-�  �BM&/       malorum     p���fU  0���fU  ��cillum dolore eu fugiat nulla pariatur olupate velit esse U  ��˝-�  �BM&/       malorum     ����fU  P���fU  Ќ�cillum dolore eu fugiat nulla pariatur olupate velit esse U  ��˝-�  �BM&/       malorum     @���fU  ����fU  ���cillum dolore eu fugiat nulla pariatur olupate velit esse U  ��g�-�  ejM&/       Workout     0���fU  ����fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��g�-�  ejM&/       Workout     ���fU  ����fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��g�-�  ejM&/       Workout     ����fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��g�-�  ejM&/       Workout     ����fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��-�  d�M&/      Meeting     P���fU  ���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  P���fU  ���fU  P��-�  �M&/       bonorum                        Excepteur sint occaecat cupidatat non proident               P��-�  �M&/       bonorum     �7��fU  `8��fU   9�Excepteur sint occaecat cupidatat non proident ��fU  P>��fU  P��-�  �M&/       bonorum     :��fU  �:��fU  ;�Excepteur sint occaecat cupidatat non proident ��fU  �>��fU  P��-�  �M&/       bonorum     p|��fU  0}��fU  �}�Excepteur sint occaecat cupidatat non proident ��fU  ����fU  \�)�-�  ��M&/      bonorum     �&��fU  p'��fU  �)�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   D�Π-�  �N&/      Appointment ���fU  P ��fU  �"�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   rp�-�  D1N&/      Birthday    0���fU  ����fU  0��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ,"�-�  m[N&/      Meeting     @f��fU   g��fU  �j�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �鐢-�  {N&/      exercitation                   Excepteur sint occaecat cupidatat non proident                "£-�  @�N&/       bonorum     ����fU  ����fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  "£-�  @�N&/       bonorum     z��fU  �z��fU  {�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �_�-�  �O&/      bonorum     �`��fU  @a��fU  �a�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ����-�  c@O&/       Appointment ����fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ����-�  c@O&/       Appointment  ���fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   t=5�-�  �iO&/      malorum     ����fU  ����fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq    �˦-�  `�O&/       Workout fU  ����fU  ����fU  @��Excepteur sint occaecat cupidatat non proident ��fU  `���fU  �˦-�  `�O&/       Workout     _��fU  �_��fU  �`�Excepteur sint occaecat cupidatat non proident ��fU  e��fU  �˦-�  `�O&/       Workout fU   ���fU  ����fU   ��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  �˦-�  `�O&/       Workout      f��fU  �f��fU  �g�Excepteur sint occaecat cupidatat non proident ��fU  `w��fU  )Oئ-�  ��O&/       Birthday    �L��fU  �M��fU  pN�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  +Oئ-�  ��O&/       Birthday    ����fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat iq   -Oئ-�  ��O&/       Birthday    ����fU   ���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat iq   /Oئ-�  ��O&/       Birthday    �T��fU  0���fU   V�ullamco laboris nisi ut aliquip ex ea commodo consequat iq   ��p�-�  ��O&/      exercitation ��fU   ��fU  ��cillum dolore eu fugiat nulla pariatur ��fU   ��fU  �!��fU  �-�  ��O&/      malorum     `��fU  ���fU  ��cillum dolore eu fugiat nulla pariatur ��fU  ���fU  0 ��fU  �0�-�  ��O&/       Appointment P���fU  ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �0�-�  ��O&/       Appointment �C��fU  @D��fU   E�Duis aute irure dolor in rehendert in volupate velit esse U  �0�-�  ��O&/       Appointment �4��fU  `5��fU   6�Duis aute irure dolor in rehendert in volupate velit esse U  �0�-�  ��O&/       Appointment �P��fU  `Q��fU   R�Duis aute irure dolor in rehendert in volupate velit esse U  <q��-�  wP&/      malorum tion ���fU  ����fU  ���cillum dolore eu fugiat nulla pariatur roident onsequat �fU  ��*�-�  �+P&/       exercitation d��fU  `e��fU   f�cillum dolore eu fugiat nulla pariatur ��fU  `j��fU  �j��fU  ��*�-�  �+P&/       exercitation j��fU  �j��fU  �v�cillum dolore eu fugiat nulla pariatur et dolor magna aliq   ��*�-�  �+P&/       exercitation \��fU  �]��fU  p^�cillum dolore eu fugiat nulla pariatur et dolor magna aliq   ��*�-�  �+P&/       exercitation u��fU  �u��fU  0v�cillum dolore eu fugiat nulla pariatur et dolor magna aliq   ©-�  uRP&/       Workout                        cillum dolore eu fugiat nulla pariatur                       	©-�  uRP&/       Workout     m��fU  �m��fU  n�cillum dolore eu fugiat nulla pariatur ��fU   q��fU  �q��fU  
©-�  uRP&/       Workout     `|��fU  �|��fU  �}�cillum dolore eu fugiat nulla pariatur ��fU  ����fU  `���fU  ©-�  uRP&/       Workout     p���fU  ����fU  p��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  p���fU  ^�-�  _zP&/       Appointment                    sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ^�-�  _zP&/       Appointment ����fU  ����fU  0��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ^�-�  _zP&/       Appointment 0J��fU  �J��fU  0K�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ^�-�  _zP&/       Appointment ����fU  `���fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   L�-�  �P&/      Meeting     ����fU  p���fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  oD��-�  U�P&/      Meeting     �?��fU   @��fU  �@�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ���-�  �P&/       consectetur ����fU  `���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  ���-�  �P&/       consectetur P���fU  ���fU  п�sunt in culpa qui offici desunt molit aim id est laborum. U  ���-�  �P&/       consectetur ���fU  ����fU  p��sunt in culpa qui offici desunt molit aim id est laborum. U  ���-�  �P&/       consectetur ����fU  `���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  ���-�  ~�P&/      bonorum     ���fU  P��fU  �sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �k�-�  j�[&/       Appointment 0��fU  ���fU  �	�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �k�-�  j�[&/       Appointment ���fU  ����fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �k�-�  j�[&/       Appointment  ��fU  ���fU  `�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �k�-�  j�[&/       Appointment @���fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �$x�-�  ��[&/       bonorum     :��fU  �:��fU  ;�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �$x�-�  ��[&/       bonorum     ����fU  `���fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �|�-�  ��[&/      exercitation ���fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  в��-�  ��[&/       Workout fU   ���fU  ����fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Ҳ��-�  ��[&/       Workout                        sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Բ��-�  ��[&/       Workout     ���fU  ����fU  0��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ز��-�  ��[&/       Workout     �y��fU   z��fU  �z�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �y�-�  ��[&/      bonorum     0T��fU  �T��fU  pU�Excepteur sint occaecat cupidatat non proident ��fU  �Z��fU  侞�-�  \&/      Workout     p���fU  0���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU  p���fU  �/�-�  95\&/      bonorum     `���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ��i�-�  ��\&/       Appointment p���fU  0���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��i�-�  ��\&/       Appointment л��fU  ����fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��i�-�  ��\&/       Appointment  ���fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��i�-�  ��\&/       Appointment �|��fU   }��fU  �}�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  $Em�-�  x�\&/      consectetur @��fU   ��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ����-�  �\&/       Birthday    @���fU   ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  �	��fU  ����-�  �\&/       Birthday    pN��fU  0O��fU  �O�Excepteur sint occaecat cupidatat non proident ��fU  �T��fU  ����-�  �\&/       Birthday    0K��fU  �K��fU  0L�Excepteur sint occaecat cupidatat non proident ��fU  PO��fU  ����-�  �\&/       Birthday    p���fU  0���fU  ��Excepteur sint occaecat cupidatat non proident ��fU  p���fU  ��-�   �\&/       bonorum     @���fU   ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  �	��fU  ��-�   �\&/       bonorum     ����fU   ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  `���fU  ��-�   �\&/       bonorum     ����fU   ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  @���fU  ��-�   �\&/       bonorum     ���fU  `��fU  ��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  �*�-�  >�\&/      malorum fU  @���fU  ���fU  p��sunt in culpa qui offici desunt molit aim id est laborum. U  ��K�-�  � ]&/       exercitation                   sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��K�-�  � ]&/       exercitation ���fU  ����fU  p��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��K�-�  � ]&/       exercitation ���fU  ����fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��K�-�  � ]&/       exercitation ���fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   L3��-�  a#]&/      Birthday U  �}��fU  �~��fU  p�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  kpd�-�  �H]&/       Meeting ent Pg��fU  �g��fU  Ph�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  mpd�-�  �H]&/       Meeting ent ���fU   	��fU  �	�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  x�s�-�  �L]&/       Birthday    ���fU  P��fU  �cillum dolore eu fugiat nulla pariatur ��fU  0��fU  ���fU  y�s�-�  �L]&/       Birthday ion ���fU  ����fU  ���cillum dolore eu fugiat nulla pariatur olupate velit esse U  z�s�-�  �L]&/       Birthday ion ���fU  О��fU  ���cillum dolore eu fugiat nulla pariatur olupate velit esse U  |�s�-�  �L]&/       Birthday ion                   cillum dolore eu fugiat nulla pariatur olupate velit esse    ���-�  ��]&/      Birthday    �N��fU  PO��fU  �O�Excepteur sint occaecat cupidatat non proident ��fU  �S��fU  K%�-�  ��]&/      Workout fU  ����fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  $��-�  �]&/      Workout fU  @��fU   ��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   )(��-�  )�]&/       Meeting     �E��fU  `F��fU  �F�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  *(��-�  )�]&/       Meeting     �<��fU   =��fU  �=�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  1i�-�  �^&/       Birthday ur  ��fU  ���fU   �sunt in culpa qui offici desunt molit aim id est laborum. U  2i�-�  �^&/       Birthday ur  ���fU  ����fU   ��sunt in culpa qui offici desunt molit aim id est laborum. U  ��v�-�  ^&/      bonorum fU  ����fU  p���fU  P��Duis aute irure dolor in rehendert in volupate velit esse U  P���-�  �W^&/       Birthday    ����fU  p���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  0���fU  ����fU  Q���-�  �W^&/       Birthday    @���fU  ����fU  @��cillum dolore eu fugiat nulla pariatur ommodo consequat . U  <T%�-�  W�^&/      consectetur `|��fU  �|��fU  �}�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Ec��-�  ��^&/      bonorum     @���fU   ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU   ��-�  �^&/       exercitation ���fU  p���fU  P��cillum dolore eu fugiat nulla pariatur ��fU  P���fU  ���fU   ��-�  �^&/       exercitation ���fU  ����fU  ���cillum dolore eu fugiat nulla pariatur ��fU  `���fU   ���fU   ��-�  �^&/       exercitation ���fU  ����fU  ���cillum dolore eu fugiat nulla pariatur ��fU  `���fU   ���fU   ��-�  �^&/       exercitation ��fU  `��fU  ��cillum dolore eu fugiat nulla pariatur ��fU   ��fU  ���fU  �S�-�  ��^&/       exercitation ���fU  @���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  �S�-�  ��^&/       exercitation 8��fU  �9��fU  :�sunt in culpa qui offici desunt molit aim id est laborum. U  �Bn�-�  ��^&/       Meeting ent  6��fU  �6��fU  �7�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �Bn�-�  ��^&/       Meeting ent @���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �Bn�-�  ��^&/       Meeting ent @���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �Bn�-�  ��^&/       Meeting ent ����fU  ����fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��r�-�  ��^&/       bonorum fU  ����fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��r�-�  ��^&/       bonorum     D��fU  �D��fU  �G�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��r�-�  ��^&/       bonorum     ���fU  ���fU  p�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU   �r�-�  ��^&/       bonorum      R��fU  �R��fU   S�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ,#t�-�  �^&/      Appointment                    Lorem ipsum dolor sit amet, consectetur adipiscing elit      (��-�  ��^&/       exercitation 1��fU  �1��fU  �2�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  )��-�  ��^&/       exercitation 5��fU  �5��fU  P6�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  *��-�  ��^&/       exercitation ���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  +��-�  ��^&/       exercitation 7��fU  �7��fU  @8�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  $���-�  �_&/      malorum                        Lorem ipsum dolor sit amet, consectetur adipiscing elit      �J��-�  a"_&/       Appointment ���fU  P��fU  �Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �J��-�  a"_&/       Appointment �@��fU  @A��fU  �A�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �J��-�  a"_&/       Appointment P7��fU  �7��fU  �8�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �J��-�  a"_&/       Appointment p"��fU  0#��fU  �#�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ���-�  Xi_&/       Birthday    ���fU  Ћ��fU  Џ�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ���-�  Xi_&/       Birthday    ���fU  P��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ���-�  Xi_&/       Birthday     ��fU  ���fU   �ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ���-�  Xi_&/       Birthday    ����fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ㋾�-�  ,l_&/       malorum     ����fU  P���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  拾�-�  ,l_&/       malorum     ����fU  P���fU  Ќ�Duis aute irure dolor in rehendert in volupate velit esse U  P��-�  !p_&/      Birthday    ����fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �Mf�-�  �_&/      bonorum     ���fU  Ћ��fU  Џ�Duis aute irure dolor in rehendert in volupate velit esse U  l���-�  չ_&/      consectetur ���fU  Ћ��fU  Џ�Excepteur sint occaecat cupidatat non proident ��fU  0���fU  z�-�  �_&/      consectetur <��fU  �<��fU  �=�sunt in culpa qui offici desunt molit aim id est laborum. U  A��-�  ��_&/       malorum     ���fU  ����fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  B��-�  ��_&/       malorum     P���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �/�-�  	`&/      Birthday U  �s��fU  pt��fU  0u�cillum dolore eu fugiat nulla pariatur ��fU  px��fU  0y��fU  ����-�  g1`&/      Birthday U  P���fU  ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  �I�-�  =T`&/      Meeting     �O��fU  pP��fU  0Q�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   0SS�-�  �V`&/       malorum fU  ����fU  `���fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  2SS�-�  �V`&/       malorum fU  л��fU  ����fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  3SS�-�  �V`&/       malorum     ���fU  �	��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  4SS�-�  �V`&/       malorum     ����fU  `���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  ��.�  Zk&/      Workout      ���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  (�.�  �1k&/       Appointment                    ullamco laboris nisi ut aliquip ex ea commodo consequat      )�.�  �1k&/       Appointment ����fU  `���fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  *�.�  �1k&/       Appointment  R��fU  �R��fU   S�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  +�.�  �1k&/       Appointment ���fU  ����fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  Z�4.�  Qk&/      Birthday U  @���fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  �k6.�  �Qk&/       Workout fU  �n��fU  �o��fU  `p�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �k6.�  �Qk&/       Workout ent 0���fU  ����fU  `��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �k6.�  �Qk&/       Workout ent �-��fU  �.��fU  �C�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �k6.�  �Qk&/       Workout ent pU��fU  �`��fU  0W�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �mQ.�  nXk&/       malorum fU  ���fU  P��fU  �ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �mQ.�  nXk&/       malorum tur п��fU  ����fU  P��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �mQ.�  nXk&/       malorum tur  ���fU  ����fU  P��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �mQ.�  nXk&/       malorum tur @���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �K�.�  �yk&/       consectetur                    cillum dolore eu fugiat nulla pariatur                       �K�.�  �yk&/       consectetur ���fU  ����fU  P��cillum dolore eu fugiat nulla pariatur ��fU  ���fU  ����fU  �K�.�  �yk&/       consectetur �&��fU  p'��fU  �)�cillum dolore eu fugiat nulla pariatur ��fU   5��fU  �5��fU  �K�.�  �yk&/       consectetur ����fU  ����fU  0��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  `���fU  P�v.�  ��k&/       consectetur p���fU  ���fU  p��Excepteur sint occaecat cupidatat non proident ��fU  p���fU  Q�v.�  ��k&/       consectetur  0��fU  �0��fU  P1�Excepteur sint occaecat cupidatat non proident ��fU  `5��fU  �C.�  ��k&/       Birthday    @��fU   ��fU  ��Excepteur sint occaecat cupidatat non proident ��fU  �!��fU  �C.�  ��k&/       Birthday nt pN��fU  0O��fU  �O�Excepteur sint occaecat cupidatat non proident onsequat �fU  �C.�  ��k&/       Birthday nt �@��fU  PA��fU  B�Excepteur sint occaecat cupidatat non proident onsequat �fU  �C.�  ��k&/       Birthday nt P[��fU  \��fU  �\�Excepteur sint occaecat cupidatat non proident onsequat �fU  O=.�  ��k&/      exercitation ���fU  `���fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  !c�.�  4�k&/       Workout     `���fU  ����fU  `��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   "c�.�  4�k&/       Workout     �A��fU   B��fU  �B�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   p�.�  ��k&/      Appointment D��fU  �D��fU  �G�cillum dolore eu fugiat nulla pariatur ��fU  U��fU  �U��fU  P�C.�  �l&/       Appointment                    cillum dolore eu fugiat nulla pariatur                       Q�C.�  �l&/       Appointment  E��fU  �E��fU  �F�cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  R�C.�  �l&/       Appointment                    cillum dolore eu fugiat nulla pariatur ommodo consequat      T�C.�  �l&/       Appointment �A��fU   B��fU  �B�cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  �jF.�  8l&/       Birthday    �=��fU   >��fU  �>�Excepteur sint occaecat cupidatat non proident ��fU  `B��fU  �jF.�  8l&/       Birthday    0���fU  ����fU  0��Excepteur sint occaecat cupidatat non proident ��fU   ���fU  ��.�  �:l&/       bonorum fU  ����fU  0���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  ��.�  �:l&/       bonorum      '��fU  �'��fU  P(�sunt in culpa qui offici desunt molit aim id est laborum. U  \�k.�  Kel&/      bonorum fU  B��fU  pL��fU  �C�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �Wt.�  �gl&/       Workout     p���fU  0���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  �Wt.�  �gl&/       Workout  ur `���fU  ����fU  ���sunt in culpa qui offici desunt molit aim id est laborum.    �Wt.�  �gl&/       Workout  ur ����fU  0���fU  ���sunt in culpa qui offici desunt molit aim id est laborum.    �Wt.�  �gl&/       Workout  ur  ���fU  ����fU  `��sunt in culpa qui offici desunt molit aim id est laborum.    ��.�  �jl&/       consectetur `���fU  ����fU  ���Excepteur sint occaecat cupidatat non proident ��fU  `���fU  ��.�  �jl&/       consectetur `r��fU   s��fU  �s�Excepteur sint occaecat cupidatat non proident ��fU  �w��fU  ��.�  �jl&/       consectetur ����fU  ���fU  �o�Excepteur sint occaecat cupidatat non proident ��fU  pt��fU  ��.�  �jl&/       consectetur 0���fU  ����fU  0��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  ��.�  o�l&/       malorum                        Duis aute irure dolor in rehendert in volupate velit esse    ��.�  o�l&/       malorum     �*��fU  �+��fU  P,�Duis aute irure dolor in rehendert in volupate velit esse U  ��.�  o�l&/       malorum     `3��fU   4��fU  �4�Duis aute irure dolor in rehendert in volupate velit esse U  ��.�  o�l&/       malorum     �A��fU  `B��fU  �B�Duis aute irure dolor in rehendert in volupate velit esse U  t��.�  jm&/      Meeting fU  ����fU  `���fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  T�f.�  �(m&/      bonorum     ����fU  ���fU  л�Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �_�.�  -Nm&/       exercitation                   cillum dolore eu fugiat nulla pariatur                       �_�.�  -Nm&/       exercitation ���fU   ���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU   ���fU  �_�.�  -Nm&/       exercitation ���fU  ���fU  p��cillum dolore eu fugiat nulla pariatur ��fU  @���fU  ���fU  �_�.�  -Nm&/       exercitation ���fU  ���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  0���fU  ����fU  ���.�  �Om&/      Workout fU  ����fU   ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �q.�  �Pm&/       exercitation                   sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �q.�  �Pm&/       exercitation D��fU  �D��fU  �G�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �q.�  �Pm&/       exercitation  ��fU  P!��fU  �!�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �q.�  �Pm&/       exercitation ��fU  �U��fU   �sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �^�.�  tm&/       consectetur 0��fU  ���fU  �	�cillum dolore eu fugiat nulla pariatur ��fU  ���fU  ���fU  �^�.�  tm&/       consectetur ����fU  p���fU  0��cillum dolore eu fugiat nulla pariatur ��fU  ���fU  ����fU  �^�.�  tm&/       consectetur ����fU  p���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  0���fU  ����fU  �^�.�  tm&/       consectetur 0���fU  Н��fU  ���cillum dolore eu fugiat nulla pariatur ��fU  @���fU  ����fU  ��".�  P�m&/       Workout     �y��fU  pz��fU  �z�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��".�  P�m&/       Workout      R��fU  �R��fU   S�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   @ $.�  ��m&/       Meeting fU  �x��fU  py��fU  0}�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  B $.�  ��m&/       Meeting tion ���fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat . U  D $.�  ��m&/       Meeting tion 8��fU  P9��fU  �9�ullamco laboris nisi ut aliquip ex ea commodo consequat . U  G $.�  ��m&/       Meeting tion R��fU  �R��fU   S�ullamco laboris nisi ut aliquip ex ea commodo consequat . U  1L+.�  ~�m&/       Workout     ���fU  P��fU  �Excepteur sint occaecat cupidatat non proident ��fU  ���fU  3L+.�  ~�m&/       Workout fU   ���fU  ���fU  `��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  5L+.�  ~�m&/       Workout     ���fU  ����fU   ��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  8L+.�  ~�m&/       Workout     ����fU   ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  )��.�  I�m&/       malorum     `��fU   ��fU  P�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   *��.�  I�m&/       malorum tur �E��fU  pF��fU  0G�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   +��.�  I�m&/       malorum tur �?��fU  `@��fU  �@�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ,��.�  I�m&/       malorum tur �C��fU  @D��fU   E�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   $��.�  X�m&/      consectetur                    sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Q,a.�  ��m&/       malorum fU  �!��fU  P"��fU  #�Excepteur sint occaecat cupidatat non proident ��fU  �'��fU  S,a.�  ��m&/       malorum     ����fU  P���fU  ��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  U,a.�  ��m&/       malorum     P���fU  ����fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  X,a.�  ��m&/       malorum     ����fU  @���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  @���fU  �l.�  ��m&/      Birthday    `���fU   ���fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Ёr.�  B�m&/       bonorum                        Excepteur sint occaecat cupidatat non proident               ҁr.�  B�m&/       bonorum     �4��fU  `5��fU   6�Excepteur sint occaecat cupidatat non proident ��fU  �;��fU  ԁr.�  B�m&/       bonorum      ���fU  ���fU  `��Excepteur sint occaecat cupidatat non proident ��fU   ���fU  ׁr.�  B�m&/       bonorum     �~��fU  `��fU   ��Excepteur sint occaecat cupidatat non proident ��fU  `���fU  �a�.�  k8n&/       Workout fU  ����fU  ����fU  @��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �a�.�  k8n&/       Workout      ���fU  ����fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �a�.�  k8n&/       Workout     `���fU  ����fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �a�.�  k8n&/       Workout      ��fU  ���fU  P�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   � .�  :^n&/      bonorum                        Duis aute irure dolor in rehendert in volupate velit esse    1�4.�  ~cn&/       bonorum     ����fU  P���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  P��fU  2�4.�  ~cn&/       bonorum     ���fU  �	��fU  ��Excepteur sint occaecat cupidatat non proident ��fU  ��fU  X�.�  �n&/       Birthday U  ����fU  ����fU  @��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   [�.�  �n&/       Birthday    ���fU  p���fU  0��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ^�.�  �n&/       Birthday    ���fU  `��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   b�.�  �n&/       Birthday    P��fU  ���fU  P�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Z��.�  ��n&/       malorum tion ���fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ]��.�  ��n&/       malorum tion ��fU  ���fU  0�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  `��.�  ��n&/       malorum tion ��fU  ���fU   �ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  d��.�  ��n&/       malorum tion ��fU  P��fU  �ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��.�  �n&/       malorum     P��fU  ��fU  `�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��.�  �n&/       malorum     `���fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��.�  �n&/       malorum     ����fU  @���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��.�  �n&/       malorum     ���fU  ��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ɴ�.�  x�n&/       consectetur 00��fU  �0��fU  P1�cillum dolore eu fugiat nulla pariatur ��fU  P5��fU  �5��fU  ʹ�.�  x�n&/       consectetur  ���fU   ���fU   ��cillum dolore eu fugiat nulla pariatur ��fU   ���fU  ����fU  hzk .�  �n&/       bonorum fU  �+��fU  p,��fU  �,�sunt in culpa qui offici desunt molit aim id est laborum. U  izk .�  �n&/       bonorum     ����fU  ����fU  0��sunt in culpa qui offici desunt molit aim id est laborum. U  jzk .�  �n&/       bonorum     @��fU   ��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  kzk .�  �n&/       bonorum fU  ����fU  `���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  ��!.�  ��n&/       Workout fU  `���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��!.�  ��n&/       Workout     ����fU  p���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��!.�  ��n&/       Workout     �~��fU  P��fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��!.�  ��n&/       Workout fU  �N��fU   O��fU  �O�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �:�!.�   o&/       Birthday    ����fU   ���fU  P��cillum dolore eu fugiat nulla pariatur ��fU  л��fU  ����fU  �:�!.�   o&/       Birthday ur p���fU  0���fU  ��cillum dolore eu fugiat nulla pariatur im id est laborum. U  �:�!.�   o&/       Birthday ur ����fU  p���fU  0��cillum dolore eu fugiat nulla pariatur im id est laborum. U  �:�!.�   o&/       Birthday ur `���fU  ���fU  `��cillum dolore eu fugiat nulla pariatur im id est laborum. U  ���!.�  so&/      exercitation J��fU  �K��fU  V�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   mI#.�  �no&/       Appointment ����fU  `���fU   ��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  `���fU  
mI#.�  �no&/       Appointment  ��fU  ���fU  P�cillum dolore eu fugiat nulla pariatur im id est laborum. U  %Z#.�  8so&/      Birthday    ����fU   ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  l¡M.�  Fz&/      Meeting     �&��fU  p'��fU  �)�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��N.�  ��z&/      consectetur P���fU  ���fU  п�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  |�uO.�  ߽z&/      Meeting     P��fU  ��fU  `�Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  �G�O.�  Z�z&/       bonorum     �o��fU  ����fU  Pq�Duis aute irure dolor in rehendert in volupate velit esse U  �G�O.�  Z�z&/       bonorum     ��fU  ���fU  p�Duis aute irure dolor in rehendert in volupate velit esse U  t��P.�  j
{&/      Appointment `���fU   ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  )��P.�  	{&/       exercitation #��fU  p$��fU  �$�Excepteur sint occaecat cupidatat non proident ��fU  �(��fU  *��P.�  	{&/       exercitation )��fU  *��fU  �*�Excepteur sint occaecat cupidatat non proident ��fU  @D��fU  �)9Q.�  s1{&/      Appointment P���fU  ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �8�Q.�  y\{&/       bonorum      ��fU  ���fU   �Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �8�Q.�  y\{&/       bonorum tur �"��fU  `#��fU  �#�Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  ���Q.�  /^{&/      malorum                        Duis aute irure dolor in rehendert in volupate velit esse    aR.�  5}{&/       Workout                        ullamco laboris nisi ut aliquip ex ea commodo consequat      
aR.�  5}{&/       Workout     @f��fU   g��fU  �j�ullamco laboris nisi ut aliquip ex ea commodo consequat iq   aR.�  5}{&/       Workout     �*��fU  �+��fU  P,�ullamco laboris nisi ut aliquip ex ea commodo consequat iq   aR.�  5}{&/       Workout     � ��fU  0!��fU  �!�ullamco laboris nisi ut aliquip ex ea commodo consequat iq   �NuR.�  b�{&/       exercitation ���fU  ���fU  У�Excepteur sint occaecat cupidatat non proident ��fU  P���fU  �NuR.�  b�{&/       exercitation ��fU  `��fU  ��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  �NuR.�  b�{&/       exercitation ���fU  ����fU  `��Excepteur sint occaecat cupidatat non proident ��fU  `���fU  �NuR.�  b�{&/       exercitation ���fU  P���fU  p��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  K�S.�  ��{&/       Workout     ����fU  @���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  N�S.�  ��{&/       Workout     ���fU  p���fU  0��ullamco laboris nisi ut aliquip ex ea commodo consequat e U  �`S.�  !�{&/       malorum     @f��fU   g��fU  �j�Duis aute irure dolor in rehendert in volupate velit esse U  �`S.�  !�{&/       malorum     ���fU  ����fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  �`S.�  !�{&/       malorum      ���fU  ����fU   x�Duis aute irure dolor in rehendert in volupate velit esse U  �`S.�  !�{&/       malorum fU  P���fU  Р��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  ��S.�  6�{&/       Workout     P���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��S.�  6�{&/       Workout fU  ���fU  ��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ly�S.�  u�{&/      consectetur                    ullamco laboris nisi ut aliquip ex ea commodo consequat      �6T.�  G�{&/      bonorum     �~��fU  `��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ���T.�  �|&/       Birthday    �,��fU  �-��fU  p.�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ���T.�  �|&/       Birthday nt �-��fU  p.��fU   /�Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  ���T.�  �|&/       Birthday nt P(��fU  �(��fU  P)�Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  ���T.�  �|&/       Birthday nt �'��fU  �(��fU  )�Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  ���T.�  ~ |&/      Workout                        Excepteur sint occaecat cupidatat non proident               tI�U.�  Ji|&/      Birthday U  0���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  P��V.�  ��|&/       Birthday    �C��fU  @D��fU   E�cillum dolore eu fugiat nulla pariatur ��fU  �I��fU  @J��fU  Q��V.�  ��|&/       Birthday    �6��fU  `7��fU  �7�cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  R��V.�  ��|&/       Birthday    �4��fU  `5��fU  �5�cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  S��V.�  ��|&/       Birthday    01��fU  �1��fU  `2�cillum dolore eu fugiat nulla pariatur ommodo consequat �fU  T�3W.�  V�|&/      Meeting                        sunt in culpa qui offici desunt molit aim id est laborum.    D�W.�  l�|&/      Meeting     �,��fU  @-��fU  �-�cillum dolore eu fugiat nulla pariatur ��fU  P1��fU  �1��fU  y"�W.�  ��|&/       Birthday    ���fU  p���fU  ��cillum dolore eu fugiat nulla pariatur ��fU  @���fU  ����fU  z"�W.�  ��|&/       Birthday    �,��fU  P-��fU  �-�cillum dolore eu fugiat nulla pariatur et dolor magna aliq   |k�X.�  _+}&/      Appointment �n��fU  �o��fU  `p�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  وY.�  #R}&/      Appointment                    cillum dolore eu fugiat nulla pariatur                       ��1Z.�  m}}&/       Workout fU  P���fU  ����fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��1Z.�  m}}&/       Workout fU  ����fU  ����fU  @��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��1Z.�  m}}&/       Workout     У��fU  ����fU  P��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ��1Z.�  m}}&/       Workout     ����fU  `���fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  W�BZ.�  ��}&/      Workout     ���fU  ����fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  ���Z.�  N�}&/       Birthday U  ����fU  ����fU  @��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ���Z.�  N�}&/       Birthday nt ���fU  ����fU  p��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ٓV[.�  W�}&/       Appointment                    ullamco laboris nisi ut aliquip ex ea commodo consequat      ړV[.�  W�}&/       Appointment �E��fU  �F��fU   G�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ۓV[.�  W�}&/       Appointment  ��fU  ���fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ݓV[.�  W�}&/       Appointment p��fU  0��fU   �ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ,QX[.�  ��}&/       Workout     "��fU  �"��fU  #�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   .QX[.�  ��}&/       Workout     ����fU  @���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   4�`[.�  ��}&/      consectetur                    sed do eiusmo tempo incidunt ut labore et dolor magna aliq   T�	\.�  6�}&/      malorum fU  ���fU  Ћ��fU  Џ�Excepteur sint occaecat cupidatat non proident ��fU  0���fU  �*].�  @~&/      exercitation ��fU  ��fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ,b�].�  mc~&/      Birthday U  ����fU  `���fU  ��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �].�   e~&/       Meeting     �L��fU  @M��fU   N�Duis aute irure dolor in rehendert in volupate velit esse U  
�].�   e~&/       Meeting ent ����fU  0���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �+�].�  i~&/       malorum     B��fU  pL��fU  �C�Duis aute irure dolor in rehendert in volupate velit esse U  �+�].�  i~&/       malorum     ����fU  P���fU  ���Duis aute irure dolor in rehendert in volupate velit esse    �+�].�  i~&/       malorum     P��fU  ��fU  0/�Duis aute irure dolor in rehendert in volupate velit esse    �+�].�  i~&/       malorum      ���fU  ����fU   ��Duis aute irure dolor in rehendert in volupate velit esse    Jc�].�  ]k~&/       Appointment  ���fU  ����fU  `��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  Lc�].�  ]k~&/       Appointment 0��fU  ���fU  0�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  Nc�].�  ]k~&/       Appointment ���fU  ����fU  ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  Qc�].�  ]k~&/       Appointment ����fU  ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU   �^.�  Է~&/       consectetur ����fU  @���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  !�^.�  Է~&/       consectetur �O��fU  PP��fU  �P�sunt in culpa qui offici desunt molit aim id est laborum. U  ��t�.�  D؉&/       exercitation ��fU  P��fU   �sunt in culpa qui offici desunt molit aim id est laborum. U  ��t�.�  D؉&/       exercitation 
��fU  �
��fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  H0�.�  }��&/       exercitation                   Excepteur sint occaecat cupidatat non proident               I0�.�  }��&/       exercitation ���fU  p���fU  0��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  J0�.�  }��&/       exercitation ���fU  ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  K0�.�  }��&/       exercitation ���fU  Н��fU  P��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  H���.�  �)�&/       Birthday     ���fU  ����fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  K���.�  �)�&/       Birthday    ���fU  ���fU  `�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �o��.�  Z*�&/       malorum     �O��fU  pP��fU  0Q�Duis aute irure dolor in rehendert in volupate velit esse U  �o��.�  Z*�&/       malorum     ����fU  P���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  F-��.�  �*�&/      exercitation A��fU  @B��fU  �B�Duis aute irure dolor in rehendert in volupate velit esse U  IE;�.�  �L�&/       Meeting tur z��fU  �z��fU  {�Duis aute irure dolor in rehendert in volupate velit esse U  JE;�.�  �L�&/       Meeting tur Ph��fU  �h��fU  �i�Duis aute irure dolor in rehendert in volupate velit esse U  \LC�.�  �N�&/      consectetur                    Lorem ipsum dolor sit amet, consectetur adipiscing elit      �o،.�  �t�&/       consectetur                    Duis aute irure dolor in rehendert in volupate velit esse    �o،.�  �t�&/       consectetur Pc��fU  �c��fU  �d�Duis aute irure dolor in rehendert in volupate velit esse U  �o،.�  �t�&/       consectetur `p��fU   q��fU  �q�Duis aute irure dolor in rehendert in volupate velit esse U  �o،.�  �t�&/       consectetur @x��fU  �x��fU  �y�Duis aute irure dolor in rehendert in volupate velit esse U  �xt�.�  ˜�&/       bonorum     p^��fU  0_��fU  �_�Duis aute irure dolor in rehendert in volupate velit esse U  �xt�.�  ˜�&/       bonorum     ����fU  ����fU  `��Duis aute irure dolor in rehendert in volupate velit esse U  �xt�.�  ˜�&/       bonorum     P��fU   ��fU  P�Duis aute irure dolor in rehendert in volupate velit esse U  �xt�.�  ˜�&/       bonorum     0���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �t�.�  ~Ŋ&/      Workout     p���fU  0���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  �ñ�.�  �&/       consectetur ����fU  `���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �ñ�.�  �&/       consectetur  ��fU  ���fU   �Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �&2�.�  ��&/       Meeting                        ullamco laboris nisi ut aliquip ex ea commodo consequat      �&2�.�  ��&/       Meeting     0W��fU  �W��fU  �X�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �&2�.�  ��&/       Meeting     ����fU  P���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �&2�.�  ��&/       Meeting fU   ���fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �?�.�  n�&/      bonorum     U��fU  �U��fU  Y�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��ޏ.�  ;�&/       exercitation ���fU  ����fU  0��Duis aute irure dolor in rehendert in volupate velit esse U  ��ޏ.�  ;�&/       exercitation ���fU  ���fU  p��Duis aute irure dolor in rehendert in volupate velit esse    ���.�  g��&/      bonorum     ����fU   ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU   ��.�  ���&/       exercitation                   sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��.�  ���&/       exercitation ���fU  ����fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��.�  ���&/       exercitation ���fU  ����fU  @��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ��.�  ���&/       exercitation ���fU  ����fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   _��.�  9��&/      bonorum     �\��fU  ]��fU  �]�Excepteur sint occaecat cupidatat non proident ��fU  @a��fU  ��@�.�  G׋&/      bonorum tion ���fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �4ǒ.�  ���&/      Workout                        Excepteur sint occaecat cupidatat non proident               ��!�.�  㓌&/       Workout     ���fU  Ћ��fU  Џ�Duis aute irure dolor in rehendert in volupate velit esse U  ��!�.�  㓌&/       Workout     �D��fU  @E��fU  �E�Duis aute irure dolor in rehendert in volupate velit esse U  ��!�.�  㓌&/       Workout     P���fU  ���fU  п�Duis aute irure dolor in rehendert in volupate velit esse U  ��!�.�  㓌&/       Workout     @���fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  %�"�.�  8��&/      exercitation ���fU  ����fU  @��sunt in culpa qui offici desunt molit aim id est laborum. U  l���.�  2�&/      Birthday U  P���fU  ���fU  ���cillum dolore eu fugiat nulla pariatur ��fU  ����fU  P���fU  9���.�  �8�&/       bonorum fU  �9��fU  P:��fU  �1�Excepteur sint occaecat cupidatat non proident ��fU  �6��fU  :���.�  �8�&/       bonorum     ����fU   ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  ;���.�  �8�&/       bonorum     P��fU  ���fU  � �Excepteur sint occaecat cupidatat non proident ��fU  �$��fU  <���.�  �8�&/       bonorum     �J��fU  �K��fU  V�Excepteur sint occaecat cupidatat non proident ��fU  pP��fU  �k<�.�  W_�&/       Appointment                    ullamco laboris nisi ut aliquip ex ea commodo consequat      �k<�.�  W_�&/       Appointment                    ullamco laboris nisi ut aliquip ex ea commodo consequat e    �k<�.�  W_�&/       Appointment �x��fU  `y��fU  z�ullamco laboris nisi ut aliquip ex ea commodo consequat e    �k<�.�  W_�&/       Appointment 0���fU  ����fU  0��ullamco laboris nisi ut aliquip ex ea commodo consequat e    �TƘ.�  ���&/       bonorum     P���fU  ���fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �TƘ.�  ���&/       bonorum     `���fU   ���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �TƘ.�  ���&/       bonorum      ���fU  ����fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �TƘ.�  ���&/       bonorum     �	��fU  p
��fU   �ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��Ș.�  E��&/       malorum     @���fU   ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  �	��fU  ��Ș.�  E��&/       malorum     ���fU  P��fU  �Excepteur sint occaecat cupidatat non proident ��fU  ��fU  ��Ș.�  E��&/       malorum     �}��fU  �~��fU  p�Excepteur sint occaecat cupidatat non proident ��fU  ����fU  ��Ș.�  E��&/       malorum     0���fU  ����fU  0��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  C*Ϙ.�  脍&/       Appointment ����fU  ����fU  @��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   F*Ϙ.�  脍&/       Appointment  W��fU  �W��fU  `X�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   I*Ϙ.�  脍&/       Appointment                    sed do eiusmo tempo incidunt ut labore et dolor magna aliq   L*Ϙ.�  脍&/       Appointment  ���fU  ����fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �Ԙ.�  )��&/      consectetur p���fU  0���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  p���fU  �\�.�  ���&/       exercitation 
��fU  �
��fU  0�sunt in culpa qui offici desunt molit aim id est laborum. U  �\�.�  ���&/       exercitation ���fU   ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  !:f�.�  ���&/       Appointment @7��fU  �7��fU  p8�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  #:f�.�  ���&/       Appointment �|��fU  `}��fU  �}�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ʀ�.�  ��&/       consectetur ����fU  ����fU  @��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ʀ�.�  ��&/       consectetur  ��fU  ���fU  ��ullamco laboris nisi ut aliquip ex ea commodo consequat . U  ʀ�.�  ��&/       consectetur  s��fU  pt��fU  0u�ullamco laboris nisi ut aliquip ex ea commodo consequat . U  ʀ�.�  ��&/       consectetur  ���fU  ����fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat . U  �섚.�  ��&/       Birthday    0.��fU  �.��fU  `/�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �섚.�  ��&/       Birthday    t��fU  �t��fU  u�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   @��.�  ���&/       bonorum     p���fU  0���fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  @��.�  ���&/       bonorum ent ����fU  p���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  aP��.�  ���&/       consectetur �X��fU  pY��fU  0Z�Excepteur sint occaecat cupidatat non proident ��fU  0_��fU  cP��.�  ���&/       consectetur `��fU   ��fU  ��Excepteur sint occaecat cupidatat non proident ��fU  0#��fU  eP��.�  ���&/       consectetur �#��fU  p$��fU  �$�Excepteur sint occaecat cupidatat non proident ��fU  �(��fU  jP��.�  ���&/       consectetur �i��fU  j��fU  �j�Excepteur sint occaecat cupidatat non proident ��fU  �n��fU  B���.�  ��&/      exercitation Q��fU  �Q��fU  U�Duis aute irure dolor in rehendert in volupate velit esse U  ��&�.�  p�&/      Birthday                       cillum dolore eu fugiat nulla pariatur                       y���.�  �͘&/       Meeting     `|��fU  �|��fU  �}�sunt in culpa qui offici desunt molit aim id est laborum. U  z���.�  �͘&/       Meeting tion ���fU  ����fU  ��sunt in culpa qui offici desunt molit aim id est laborum.    
��.�  �ј&/      Appointment �R��fU  pS��fU  0T�Duis aute irure dolor in rehendert in volupate velit esse U  ,e�.�  I�&/       Workout     �A��fU  PB��fU  �B�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  .e�.�  I�&/       Workout tur �8��fU  �9��fU  :�Lorem ipsum dolor sit amet, consectetur adipiscing elit e U  	��.�  u�&/       Birthday    �L��fU  �M��fU  pN�Excepteur sint occaecat cupidatat non proident ��fU  pS��fU  
��.�  u�&/       Birthday    ���fU  Ћ��fU  Џ�Excepteur sint occaecat cupidatat non proident ��fU  0���fU  ��.�  u�&/       Birthday     ���fU  ����fU  0��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  ��.�  u�&/       Birthday    ����fU   ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  $�!�.�  8�&/      exercitation ���fU  ����fU  `��Duis aute irure dolor in rehendert in volupate velit esse U  ��5�.�  �e�&/       Birthday     ���fU  ����fU  ���cillum dolore eu fugiat nulla pariatur ��fU  `���fU   ���fU  ��5�.�  �e�&/       Birthday    @���fU  ����fU  @��cillum dolore eu fugiat nulla pariatur ��fU   ���fU  ����fU  �D�.�  ~i�&/      Appointment P��fU  ��fU  `�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ���.�  ��&/      Birthday U  P���fU  ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  P���fU  ��d�.�  T��&/      Meeting      ���fU  ����fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  A��.�  h��&/       Workout     ��fU  ���fU  p�Duis aute irure dolor in rehendert in volupate velit esse U  B��.�  h��&/       Workout     �$��fU  p%��fU  �%�Duis aute irure dolor in rehendert in volupate velit esse U  C��.�  h��&/       Workout     ���fU  @��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  D��.�  h��&/       Workout     ���fU  0��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  �$	�.�  zݙ&/      Workout                        Excepteur sint occaecat cupidatat non proident               9,��.�  S�&/       bonorum     ���fU  `���fU   ��Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  :,��.�  S�&/       bonorum tion ���fU  P���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit . U  4H��.�  �&/      Birthday                       Excepteur sint occaecat cupidatat non proident               /�D�.�  M.�&/      consectetur P��fU  ���fU  P�cillum dolore eu fugiat nulla pariatur ��fU  ���fU   ��fU  �bL�.�  :0�&/       Meeting fU  ����fU  ����fU  @��Excepteur sint occaecat cupidatat non proident ��fU  `���fU  �bL�.�  :0�&/       Meeting     n��fU  �n��fU  ���Excepteur sint occaecat cupidatat non proident ��fU   s��fU  �bL�.�  :0�&/       Meeting     `���fU  ����fU  `��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  �bL�.�  :0�&/       Meeting     ����fU  ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  �n��.�  =P�&/      Meeting     P���fU  ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   /j�.�  dy�&/      bonorum fU  ����fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  ��n�.�  �z�&/       consectetur ����fU  `���fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  ��n�.�  �z�&/       consectetur ���fU  �	��fU  ��Duis aute irure dolor in rehendert in volupate velit esse U  ��n�.�  �z�&/       consectetur ���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ��n�.�  �z�&/       consectetur �8��fU  P9��fU  �9�Duis aute irure dolor in rehendert in volupate velit esse U  ����.�  p��&/      consectetur                    Excepteur sint occaecat cupidatat non proident               � 
�.�  N��&/       exercitation                   cillum dolore eu fugiat nulla pariatur                       � 
�.�  N��&/       exercitation ���fU   ���fU  ��cillum dolore eu fugiat nulla pariatur  adipiscing elit �fU  � 
�.�  N��&/       exercitation ���fU  ����fU  ��cillum dolore eu fugiat nulla pariatur  adipiscing elit �fU  � 
�.�  N��&/       exercitation ���fU  p���fU  ��cillum dolore eu fugiat nulla pariatur  adipiscing elit �fU  |Z��.�  �ƚ&/      Appointment @���fU   ���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  ��E�.�  &�&/      Workout     B��fU  pL��fU  �C�Lorem ipsum dolor sit amet, consectetur adipiscing elit iq   0���.�  ^�&/       exercitation S��fU  �S��fU   T�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  1���.�  ^�&/       exercitation ���fU  ����fU  P��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  h�j�.�  1>�&/       malorum     0u��fU  �u��fU  0v�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   i�j�.�  1>�&/       malorum fU  ����fU  ����fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �S�.�  h�&/      malorum     p���fU  0���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ����.�  ���&/      exercitation ��fU  ���fU  p�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  ,���.�  �ܛ&/      consectetur �\��fU  �^��fU  b�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �x�.�  '�&/      malorum     `���fU  ���fU  `��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  ���fU  p��.�  f%�&/       bonorum                        sunt in culpa qui offici desunt molit aim id est laborum.    q��.�  f%�&/       bonorum fU   ���fU  ���fU  `��sunt in culpa qui offici desunt molit aim id est laborum. U  r��.�  f%�&/       bonorum     ����fU   ���fU  P��sunt in culpa qui offici desunt molit aim id est laborum. U  s��.�  f%�&/       bonorum     ����fU  @���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  ��.�  �O�&/      malorum     @���fU  ����fU  @��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  ����.�  h��&/      Meeting     `���fU  ����fU  `��sunt in culpa qui offici desunt molit aim id est laborum. U  `��.�  \��&/       Appointment ���fU  �	��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   a��.�  \��&/       Appointment 0���fU  ����fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   b��.�  \��&/       Appointment �_��fU  �k��fU  �a�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   d��.�  \��&/       Appointment `���fU  P���fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �9X�.�  �&/      Birthday                       Excepteur sint occaecat cupidatat non proident  magna aliq   qij�.�  Fǜ&/       Birthday    ����fU  p���fU  P��cillum dolore eu fugiat nulla pariatur ��fU  P���fU  ���fU  rij�.�  Fǜ&/       Birthday nt �t��fU  �u��fU   ��cillum dolore eu fugiat nulla pariatur ��fU  �z��fU  �{��fU  sij�.�  Fǜ&/       Birthday nt Pm��fU  �m��fU  Pn�cillum dolore eu fugiat nulla pariatur ��fU  Pr��fU  �r��fU  tij�.�  Fǜ&/       Birthday nt л��fU  ����fU  ��cillum dolore eu fugiat nulla pariatur ��fU  P���fU  ����fU  Y���.�  ��&/       consectetur  `��fU  Pa��fU  b�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   Z���.�  ��&/       consectetur  U��fU  �U��fU  0V�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   <�.�  W�&/      Meeting     @f��fU   g��fU  �j�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �՗�.�  p�&/      bonorum     �\��fU  �^��fU  b�Excepteur sint occaecat cupidatat non proident ��fU  �o��fU  ��1�.�  �;�&/      Appointment �&��fU  p'��fU  �)�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ��2�.�  <�&/       exercitation ���fU  ����fU  P��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  ��2�.�  <�&/       exercitation ���fU  ����fU   ��Excepteur sint occaecat cupidatat non proident ��fU  ����fU  ��2�.�  <�&/       exercitation ���fU  ����fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  ��2�.�  <�&/       exercitation ���fU   ���fU  ���Excepteur sint occaecat cupidatat non proident ��fU  ����fU  d�t /�  |�&/       consectetur P���fU  О��fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  f�t /�  |�&/       consectetur `���fU  ����fU  `��sunt in culpa qui offici desunt molit aim id est laborum. U  \�t /�  ��&/      Birthday    ����fU  ����fU   ��sunt in culpa qui offici desunt molit aim id est laborum. U  ��w /�  E�&/       Workout fU  ����fU  p���fU  0��Duis aute irure dolor in rehendert in volupate velit esse U  ��w /�  E�&/       Workout     Pn��fU   o��fU  �o�Duis aute irure dolor in rehendert in volupate velit esse U  ��w /�  E�&/       Workout     l��fU  �l��fU  m�Duis aute irure dolor in rehendert in volupate velit esse U  ��w /�  E�&/       Workout     `j��fU  �j��fU  �v�Duis aute irure dolor in rehendert in volupate velit esse U  �/�  G5�&/      Birthday                       sed do eiusmo tempo incidunt ut labore et dolor magna aliq   A�'/�  H;�&/       Appointment ����fU  `���fU  ��Duis aute irure dolor in rehendert in volupate velit esse    B�'/�  H;�&/       Appointment �y��fU   z��fU  �z�Duis aute irure dolor in rehendert in volupate velit esse    C�'/�  H;�&/       Appointment l��fU  �l��fU  `m�Duis aute irure dolor in rehendert in volupate velit esse    D�'/�  H;�&/       Appointment �}��fU   ~��fU  �~�Duis aute irure dolor in rehendert in volupate velit esse    �̜/�  KY�&/       Birthday                       Excepteur sint occaecat cupidatat non proident               �̜/�  KY�&/       Birthday    ����fU  P���fU  ���Excepteur sint occaecat cupidatat non proident  magna aliq   �̜/�  KY�&/       Birthday    �,��fU  @-��fU  �-�Excepteur sint occaecat cupidatat non proident  magna aliq   �̜/�  KY�&/       Birthday    �9��fU  p:��fU   =�Excepteur sint occaecat cupidatat non proident  magna aliq   �9/�  n��&/      bonorum     �E��fU  `F��fU  �F�Duis aute irure dolor in rehendert in volupate velit esse U   ��/�  ԧ�&/       malorum     <��fU  �<��fU  �=�ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  !��/�  ԧ�&/       malorum     `���fU  ����fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  "��/�  ԧ�&/       malorum     ����fU  ����fU   ��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  $��/�  ԧ�&/       malorum     P���fU  ���fU  p��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ���/�  s��&/      malorum     �\��fU  ]��fU  �]�Excepteur sint occaecat cupidatat non proident ��fU  @a��fU  �q/�  )Ѩ&/      malorum     ����fU  �	��fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �/�  ���&/       consectetur ����fU  P���fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  �/�  ���&/       consectetur  ���fU  н��fU  P��sunt in culpa qui offici desunt molit aim id est laborum.    �/�  ���&/       consectetur  ���fU  ����fU   ��sunt in culpa qui offici desunt molit aim id est laborum.    �/�  ���&/       consectetur  ��fU   ��fU  P�sunt in culpa qui offici desunt molit aim id est laborum.    U�/�  !��&/      Birthday    ���fU  ����fU  P��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �/�  `��&/       malorum     `j��fU  �j��fU  �v�Duis aute irure dolor in rehendert in volupate velit esse U  �/�  `��&/       malorum tion N��fU  �N��fU  �O�Duis aute irure dolor in rehendert in volupate velit esse U  �/�  `��&/       malorum tion M��fU  PN��fU  �N�Duis aute irure dolor in rehendert in volupate velit esse U  �/�  `��&/       malorum tion ��fU  ���fU  P�Duis aute irure dolor in rehendert in volupate velit esse U  ��!/�  l��&/       Meeting      x��fU  �x��fU  �y�Excepteur sint occaecat cupidatat non proident ��fU  `~��fU  ��!/�  l��&/       Meeting fU  �-��fU  p.��fU   /�Excepteur sint occaecat cupidatat non proident velit esse U  ��!/�  l��&/       Meeting      ���fU  ����fU   x�Excepteur sint occaecat cupidatat non proident velit esse U  ��!/�  l��&/       Meeting      S��fU  �S��fU   T�Excepteur sint occaecat cupidatat non proident velit esse U  h�/�  ��&/       Meeting      5��fU  �5��fU  �9�Duis aute irure dolor in rehendert in volupate velit esse U  i�/�  ��&/       Meeting  U  Ѐ��fU  P���fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  j�/�  ��&/       Meeting     ����fU  0���fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  k�/�  ��&/       Meeting     `���fU  ����fU  ���Duis aute irure dolor in rehendert in volupate velit esse U  $y�/�  �n�&/      Workout     ����fU  ����fU  `��sunt in culpa qui offici desunt molit aim id est laborum. U  ��b/�  +��&/       malorum     �'��fU  �(��fU  )�Duis aute irure dolor in rehendert in volupate velit esse U  ��b/�  +��&/       malorum      ���fU  ����fU   ��Duis aute irure dolor in rehendert in volupate velit esse U  A'n/�  ��&/       consectetur  9��fU  @C��fU  �:�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   B'n/�  ��&/       consectetur ���fU  ���fU   �sed do eiusmo tempo incidunt ut labore et dolor magna aliq   C'n/�  ��&/       consectetur 0T��fU  �T��fU  pU�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   E'n/�  ��&/       consectetur �8��fU  `9��fU   :�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �p�/�  {��&/      malorum                        sed do eiusmo tempo incidunt ut labore et dolor magna aliq   p /�  ���&/       exercitation H��fU  �H��fU  �I�sunt in culpa qui offici desunt molit aim id est laborum. U  q /�  ���&/       exercitation ���fU  ����fU  @��sunt in culpa qui offici desunt molit aim id est laborum. U  r /�  ���&/       exercitation ���fU  ���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  s /�  ���&/       exercitation ���fU  ����fU   ��sunt in culpa qui offici desunt molit aim id est laborum. U  �=�/�  �&/       bonorum     ����fU  ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �=�/�  �&/       bonorum     `���fU  ���fU  `��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �Z�/�  ��&/       Workout      ��fU  ���fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  �Z�/�  ��&/       Workout      ��fU  ���fU   �sunt in culpa qui offici desunt molit aim id est laborum.    �Z�/�  ��&/       Workout     �=��fU  P>��fU  ?�sunt in culpa qui offici desunt molit aim id est laborum.    �Z�/�  ��&/       Workout     �&��fU  `'��fU  �'�sunt in culpa qui offici desunt molit aim id est laborum.    �C�/�  �/�&/      consectetur P(��fU  �(��fU  P)�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  @O�	/�  ~�&/       consectetur                    Excepteur sint occaecat cupidatat non proident               BO�	/�  ~�&/       consectetur p��fU   ��fU  @�Excepteur sint occaecat cupidatat non proident ��fU  @��fU  CO�	/�  ~�&/       consectetur ����fU  p���fU  0��Excepteur sint occaecat cupidatat non proident ��fU  ���fU  EO�	/�  ~�&/       consectetur �d��fU  0e��fU  �e�Excepteur sint occaecat cupidatat non proident ��fU  �i��fU  =�	/�  7~�&/      Workout fU   6��fU  �6��fU  �7�sunt in culpa qui offici desunt molit aim id est laborum. U  Ē
/�  8��&/       consectetur ����fU  @���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   ƒ
/�  8��&/       consectetur ���fU  P��fU  ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �9�
/�  �&/      Meeting     ����fU  �	��fU  ���cillum dolore eu fugiat nulla pariatur ��fU   ���fU  ����fU  `ܭ
/�  |��&/       Appointment ����fU  `���fU  ���sunt in culpa qui offici desunt molit aim id est laborum. U  bܭ
/�  |��&/       Appointment  ���fU  ���fU  `��sunt in culpa qui offici desunt molit aim id est laborum.    cܭ
/�  |��&/       Appointment  ���fU  ����fU  `��sunt in culpa qui offici desunt molit aim id est laborum.    dܭ
/�  |��&/       Appointment `���fU  ���fU  `��sunt in culpa qui offici desunt molit aim id est laborum.    0{�/�  �?�&/       bonorum fU  ����fU  ����fU  @��cillum dolore eu fugiat nulla pariatur ��fU  ����fU  `���fU  2{�/�  �?�&/       bonorum     P���fU  О��fU  ���cillum dolore eu fugiat nulla pariatur ��fU  У��fU  ����fU  4{�/�  �?�&/       bonorum     P
��fU  �
��fU  ��cillum dolore eu fugiat nulla pariatur ��fU  ���fU  ��fU  6{�/�  �?�&/       bonorum      '��fU  �'��fU  P(�cillum dolore eu fugiat nulla pariatur ��fU  �+��fU  PM��fU  y,/�  �G�&/       Workout     ����fU  P���fU  ��sunt in culpa qui offici desunt molit aim id est laborum. U  {,/�  �G�&/       Workout     �*��fU  �+��fU  P,�sunt in culpa qui offici desunt molit aim id est laborum. U  },/�  �G�&/       Workout      0��fU  �0��fU  P1�sunt in culpa qui offici desunt molit aim id est laborum. U  ,/�  �G�&/       Workout     ����fU  p���fU  0��sunt in culpa qui offici desunt molit aim id est laborum. U  ���/�  6i�&/       Meeting fU  �2��fU  3��fU  �3�Excepteur sint occaecat cupidatat non proident ��fU  �7��fU  ���/�  6i�&/       Meeting     4��fU  �4��fU  P5�Excepteur sint occaecat cupidatat non proident ��fU  P9��fU  ��/�  nj�&/      exercitation ���fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   \�#/�  K��&/      Appointment �x��fU  py��fU  0}�Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �$�/�  ̵�&/       Birthday U  ����fU  ����fU  @��Duis aute irure dolor in rehendert in volupate velit esse U  �$�/�  ̵�&/       Birthday    �C��fU  @D��fU   E�Duis aute irure dolor in rehendert in volupate velit esse U  �$�/�  ̵�&/       Birthday    �B��fU  pC��fU  �C�Duis aute irure dolor in rehendert in volupate velit esse U  �$�/�  ̵�&/       Birthday    ����fU  p���fU  0��Duis aute irure dolor in rehendert in volupate velit esse U  ��/�  ּ�&/       malorum     `���fU  ���fU  `��ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  ���/�  ּ�&/       malorum     ����fU  ����fU  ���ullamco laboris nisi ut aliquip ex ea commodo consequat �fU  �r�/�  ���&/       Birthday    �^��fU  _��fU  �_�cillum dolore eu fugiat nulla pariatur ��fU   c��fU  �c��fU  �r�/�  ���&/       Birthday    ����fU  p���fU  P��cillum dolore eu fugiat nulla pariatur ��fU  P���fU  ���fU  \�s/�  K�&/      exercitation &��fU  p'��fU  �)�sunt in culpa qui offici desunt molit aim id est laborum. U  u/�  ��&/       Workout     `j��fU  �j��fU  �v�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   u/�  ��&/       Workout     ���fU  @��fU   �sed do eiusmo tempo incidunt ut labore et dolor magna aliq   u/�  ��&/       Workout     4��fU  �4��fU  P5�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   u/�  ��&/       Workout     ����fU    ��fU  � �sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �M�/�  n�&/       Birthday    P���fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �M�/�  n�&/       Birthday    ����fU   ���fU  ���sed do eiusmo tempo incidunt ut labore et dolor magna aliq   l��/�  ��&/      Appointment ����fU  `���fU   ��cillum dolore eu fugiat nulla pariatur ��fU   ���fU  ����fU  Ae�/�  ��&/       Appointment                    sunt in culpa qui offici desunt molit aim id est laborum.    Ce�/�  ��&/       Appointment �H��fU   I��fU  �I�sunt in culpa qui offici desunt molit aim id est laborum. U  xf�/�  ;0�&/       Appointment p^��fU  0_��fU  �_�Excepteur sint occaecat cupidatat non proident ��fU  `e��fU  yf�/�  ;0�&/       Appointment ����fU   ���fU  ���Excepteur sint occaecat cupidatat non proident  magna aliq   ��1/�  oV�&/      Meeting     P���fU  ���fU  ���Lorem ipsum dolor sit amet, consectetur adipiscing elit �fU  �Ƽ/�  z�&/       consectetur  ���fU  ����fU   ��sed do eiusmo tempo incidunt ut labore et dolor magna aliq   �Ƽ/�  z�&/       consectetur  K��fU  �K��fU  PL�sed do eiusmo tempo incidunt ut labore et dolor magna aliq   4	�/�  �z�&/      malorum fU  �X��fU  pY��fU  0Z�Duis aute irure dolor in rehendert in volupate velit esse U  