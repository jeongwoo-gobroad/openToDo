ps/   us/       Birthday    ���U  ���U  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   '��U  u�/   e�/       Meeting     P3 ��U  4 ��U  �7 Some_stuffs_Some_stuffs_ �U  �@ ��U  �A ��U  pE ��U  0F ��U  q�/   ��/       Birthday    `���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  У��U  4/   e/      Birthday nt `Y��U  �Y��U  �ZThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   _��U  4/   �3/       Meeting     �� ��U  p� ��U  0� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @� ��U  `_/   h_/       Some_stuffs P% ��U  & ��U  �) Some_stuffs_Some_stuffs_ �U  P3 ��U  4 ��U  �7 ��U  �8 ��U  �/   ��/      Meeting     ����U  ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��/   ��/      Some_stuffs `_ ��U   ` ��U  `d This_stuffs_This_stuffs_ �U  �n ��U  Po ��U  �t ��U  �v ��U  ��/   ��/      Appointment p���U  0 ��U  � Some_stuffs_Some_stuffs_ �U  ���U  `��U  ���U  ���U  ��/   -�/       Some_stuffs �� ��U  @ ��U   This_stuffs_This_stuffs_ �U  ���U  ���U  @��U   ��U   /   /       Birthday    � ��U  � ��U  � This_stuffs_This_stuffs_ �U  0 ��U  � ��U  � ��U  � ��U  $J/   5J/       Appointment ����U  @���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  
p/   Nq/       Workout     �� ��U  �� ��U  @� This_stuffs_This_stuffs_ �U   � ��U  �� ��U  �� ��U  @� ��U  )�/   +�/       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ��/   J�/       Meeting     p��U  ���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ��U  /   �/       Workout     ����U  p���U  ��This_stuffs_This_stuffs_ �U  ����U  ����U  0���U  ����U  �0/   �0/       Birthday     ��U  ���U  �This_stuffs_This_stuffs_ �U   ��U  ���U  �B��U  pC��U  Z/   Z/       Workout �U  ���U  ����U  0�This_stuffs_This_stuffs_ �U  p���U  ����U  ����U  0���U  ��/   ��/       Birthday nt p���U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��/   =�/       Workout     @� ��U   � ��U  �� Some_stuffs_Some_stuffs_ �U   ��U  ���U  @��U   ��U  )�/   ^�/       Some_stuffs @���U   ���U  ��justforfun_justforfun_ ��U  ����U   ���U  ����U  @���U  ��/   ��/      Meeting ffs ����U  @���U  ��justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  `���U  /   �/       Birthday    �/��U  �0��U  `1This_stuffs_This_stuffs_ �U  �3��U  �4��U   5��U  �5��U  YF/   [H/      Birthday    Ы��U  ����U  P�Some_stuffs_Some_stuffs_ �U  ���U  а��U  ����U  ���U  m/   i/       Appointment Ѕ��U  ����U  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  -�/   c�/      Some_stuffs ���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  ��/   ��/      Some_stuffs @���U  ����U  p�justforfun_justforfun_ ��U  п��U  P���U  ���U  ����U  9/   i/       Some_stuffs �8��U  @9��U  `RSome_stuffs_Some_stuffs_ �U  �<��U   =��U  �=��U  �>��U  6�#/   $�#/       Meeting     ���U  @��U  �justforfun_justforfun_ ��U  ���U  @��U  ���U  p��U  ��#/   ��#/       Birthday nt �c��U  `d��U  �dThis_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U   i��U  �$/   �$/      Workout     �Z��U   [��U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0_��U  �'$/   C,$/       Meeting �U  �h��U  0i��U  �ijustforfun_justforfun_ ��U  �k��U  `l��U  �l��U  `m��U  �W$/   �W$/      Some_stuffs P��U  ���U  �justforfun_justforfun_ ��U  ���U   ��U  � ��U  `!��U  �~$/   y$/       Birthday    �����U  `����U  ��justforfun_justforfun_ ���U  �����U  p����U  0����U  ����U  ��$/   ��$/       Some_stuffs �0��U  p1��U  �1Some_stuffs_Some_stuffs_ �U  �3��U  p4��U  �4��U  �5��U  �$/   ��$/       Appointment �� ��U  P� ��U   � This_stuffs_This_stuffs_ �U  � ��U  Ж ��U  �� ��U  p� ��U  %�$/   g�$/       Meeting     ���U  0��U  �This_stuffs_This_stuffs_ �U  `��U   ��U  ���U  `��U  5%/   9%/       Meeting     p>��U  �>��U  �?This_stuffs_This_stuffs_ �U  �t��U  `u��U  �B��U  0C��U  =%/   �<%/      Birthday    p���U  ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  h%/   !h%/       Appointment ����U  0���U  ��This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  �%/   Í%/       Meeting     �x��U  `y��U  �yjustforfun_justforfun_ ��U  �|��U  `}��U  ����U  p���U  ��%/   ��%/      Appointment �����U  @����U  ���Some_stuffs_Some_stuffs_ �U  �����U  P����U  �����U  @����U  x�%/   y�%/       Some_stuffs  ���U  ����U    justforfun_justforfun_ ��U  `��U   ��U  ���U  ���U  j &/   �&/      Workout      x��U  �x��U  �yThis_stuffs_This_stuffs_ �U   |��U  �|��U  �}��U  @~��U  x'&/   |'&/       Workout     `w��U  �w��U  �xjustforfun_justforfun_ ��U  `{��U  �{��U  �|��U  `}��U  �P&/   Q&/      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �v&/   �v&/      Some_stuffs �:��U  `;��U   <This_stuffs_This_stuffs_ �U  �?��U  `@��U   A��U  �A��U  ��&/   ��&/       Appointment ����U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��&/   ��&/       Birthday    @o��U   p��U  �pThis_stuffs_This_stuffs_ �U  �s��U  @t��U  �t��U  �u��U  ��&/   ��&/      Birthday    ���U   '��U  Pjustforfun_justforfun_ ��U  P ��U  !��U  �!��U  �"��U  j'/   �'/       Some_stuffs P����U  ����U  P��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  �7'/   �7'/      Workout      � ��U  �� ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P� ��U  h^'/   �^'/      Meeting     ���U  P��U   This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `"��U  {�'/   ��'/       Workout      N��U  �N��U  `OSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   T��U  Q�'/   )�'/      Birthday    �� ��U  p� ��U  0� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  	�'/   ��'/       Meeting ent Pg��U  �g��U  p�This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  �k��U  ��2/   '�2/       Meeting ffs  ���U  ����U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  [!3/   ["3/       Birthday    ����U  @���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �D3/   6I3/       Workout     ����U  P���U  �Some_stuffs_Some_stuffs_ �U  P���U  ���U  ����U  P���U  �m3/   �m3/       Some_stuffs �V��U  pW��U  �WThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @\��U  E�3/   ��3/       Meeting     P� ��U  @� ��U  0� This_stuffs_This_stuffs_ �U  0� ��U  �� ��U  �� ��U  p� ��U  p�3/   L�3/       Appointment @����U  ����U  P��Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ����U  F�3/   ��3/      Workout     �'��U   (��U  �(justforfun_justforfun_ ��U  �+��U  �,��U   -��U  �-��U  �4/   Z4/      Meeting     ����U  `���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  ,34/   U34/      Some_stuffs px��U  �x��U  pyjustforfun_justforfun_ ��U  p{��U  �{��U  p|��U  0}��U  �T4/   �V4/       Some_stuffs ����U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  d}4/   }4/       Meeting     P% ��U  & ��U  �) justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  �8 ��U  |�4/   ��4/       Appointment �t ��U  �v ��U  �z This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  ��4/   x�4/      Birthday    �� ��U  �� ��U   � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `� ��U  ��4/   ��4/       Workout     ����U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �5/   5/       Workout     ����U  @���U  ��Some_stuffs_Some_stuffs_ �U  ����U  @���U  ����U  @���U  }A5/   yE5/       Appointment ���U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  ag5/   m5/       Meeting ffs �����U  P����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �  ��U  ��5/   �5/       Some_stuffs � ��U  Ж ��U  �� justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  @� ��U  =�5/   �5/       Workout     ����U  p���U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��5/   �5/      Workout �U  `*��U   +��U  �+justforfun_justforfun_ ��U  �.��U  `/��U   0��U  �0��U  	6/   �6/       Meeting     �� ��U  @� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P� ��U  �06/   �06/       Some_stuffs �
��U  ���U  �"Some_stuffs_Some_stuffs_ �U   ��U  ���U   ��U  ���U  �T6/   �Q6/      Meeting     ���U  ���U  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p��U  �z6/   Zy6/       Workout     м ��U  �� ��U  P� This_stuffs_This_stuffs_ �U  P� ��U  � ��U  �� ��U  �� ��U  �6/   ۠6/       Birthday    `��U  ���U  `Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `��U  ��6/   �6/       Appointment �W��U  pX��U   YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �]��U  �6/   9�6/       Birthday    �A��U  �B��U   CThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �G��U  �7/   7/      Meeting     �t��U  �u��U   vThis_stuffs_This_stuffs_ �U   x��U  �x��U  �y��U  @z��U  �c7/   �e7/       Some_stuffs  ��U  ���U   Some_stuffs_Some_stuffs_ �U  ���U   ��U  ���U   ��U  ��7/   �7/       Appointment                    justforfun_justforfun_                                       \;B/   �;B/       Birthday    ����U  `���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �^B/   YaB/       Appointment ����U  p���U  ��This_stuffs_This_stuffs_ �U  p���U  0���U  ����U  0���U  ��B/   0�B/      Birthday U  �����U  �����U  ���Some_stuffs_Some_stuffs_ �U  �����U  @����U  �����U  @����U  4�B/   6�B/       Some_stuffs �� ��U  `� ��U   � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0� ��U  �B/   ��B/      Appointment ����U  @���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  > C/   `�B/      Workout �U  ����U  p���U   �This_stuffs_This_stuffs_ �U  P���U   ���U  ����U   ���U  p*C/   �%C/       Birthday U  �	��U  @
��U  �
Some_stuffs_Some_stuffs_ �U  ���U  @��U   ��U  ���U  hLC/   pLC/      Birthday nt �� ��U  � ��U  Ы This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  `� ��U  XpC/   hpC/      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �C/   ,�C/       Workout     `*��U   +��U  �+This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �0��U  ��C/   n�C/       Meeting      o��U  �o��U   pjustforfun_justforfun_ ��U  `r��U   s��U  �s��U  Pt��U  ��C/   ��C/       Meeting ffs ����U  0���U  ��This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ���U  �D/   �D/       Workout ent  � ��U  �� ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  -7D/   �8D/       Workout     ����U   ���U  �Some_stuffs_Some_stuffs_ �U  `���U  ���U  ����U  `���U  �bD/   &cD/      Meeting     ����U   ���U  ��Some_stuffs_Some_stuffs_ �U  ����U  ���U  ����U  0���U  ��D/   A�D/       Workout �U  ����U  ����U  `�Some_stuffs_Some_stuffs_ �U  ����U   ���U  ����U  `���U  ��D/   ۩D/       Birthday U  �����U  �����U  ���Some_stuffs_Some_stuffs_ �U  �����U  @����U  �����U  @����U  4�D/   8�D/      Some_stuffs ����U  @���U  ��This_stuffs_This_stuffs_ �U  ����U  @���U   ���U  ����U  �D/   ��D/       Workout     ���U  `��U   Some_stuffs_Some_stuffs_ �U  ���U  `��U  ���U  ���U  �#E/   �#E/       Meeting     p\��U  0]��U  �]This_stuffs_This_stuffs_ �U  �`��U  pa��U  0b��U  �b��U  /JE/   ,IE/       Meeting     0����U  �����U  P��This_stuffs_This_stuffs_ �U  �����U  �����U   ����U  �����U  ^tE/   sE/      Some_stuffs 0����U  ����U  ���This_stuffs_This_stuffs_ �U   ����U  �����U  �����U  p����U  ��E/   *�E/       Appointment `���U   ���U  ��This_stuffs_This_stuffs_ �U  ����U   ���U  ����U   ���U  �E/   |�E/       Meeting     �� ��U  P� ��U   � This_stuffs_This_stuffs_ �U  0� ��U  � ��U  �� ��U  p� ��U  ��E/   ��E/       Some_stuffs                    justforfun_justforfun_                                       
1F/   �1F/      Workout ffs P���U  П��U  ��This_stuffs_This_stuffs_ �U  ����U  0���U  ����U  0���U  �UF/   ^F/       Meeting     ����U  P���U  �Some_stuffs_Some_stuffs_ �U  ���U  Л��U  ����U  ���U  ̅F/   ޅF/       Some_stuffs  J ��U  �J ��U  �N This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ` ��U  ��F/   ��F/       Appointment �l��U  Pm��U  �mSome_stuffs_Some_stuffs_ �U  �~��U   ��U  �p��U  �q��U  �{Q/   �{Q/      Meeting     ���U  `���U   �justforfun_justforfun_ ��U  ����U  `���U  ���U  ����U  H�Q/   Y�Q/       Some_stuffs ����U  ����U  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��Q/   ��Q/       Appointment ����U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  S�Q/   ��Q/       Workout      ;��U  �;��U  �<Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   A��U  R/   xR/      Appointment  J ��U  �J ��U  �N This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ` ��U  �kR/   �hR/      Birthday    � ��U  � ��U  � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  � ��U  �R/   Q�R/      Appointment ����U  `���U  �This_stuffs_This_stuffs_ �U  ���U  б��U  ����U  ���U  ��R/   ��R/      Some_stuffs                    justforfun_justforfun_                                       �R/    �R/      Appointment � ��U  � ��U  � This_stuffs_This_stuffs_ �U   ! ��U  �! ��U  P% ��U  & ��U  S/   �S/       Meeting     ����U  P���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �(S/   �.S/      Appointment  I��U  �I��U  PJThis_stuffs_This_stuffs_ �U  pL��U  �L��U  �M��U  0N��U  1QS/   @SS/       Appointment �b��U  Pc��U  �cThis_stuffs_This_stuffs_ �U  Pf��U  �f��U  Pg��U  �g��U  ~S/   �}S/       Meeting     �. ��U  �/ ��U  P3 This_stuffs_This_stuffs_ �U  @< ��U   = ��U  �@ ��U  �A ��U  ��S/   ��S/       Appointment @���U   ���U  ��justforfun_justforfun_ ��U  p���U  ���U  ����U   ���U  ��S/   n�S/      Meeting      5��U  �5��U  �6Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `;��U  }�S/   ��S/      Some_stuffs `���U  ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  �T/   �T/       Birthday     � ��U  �� ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   � ��U  ?T/   (?T/      Meeting     о��U  P���U  ��This_stuffs_This_stuffs_ �U  @���U  ����U  ����U  @���U  `�T/   p�T/       Appointment                    justforfun_justforfun_                                       5�T/   ��T/       Meeting  fs �I��U  �J��U  `KThis_stuffs_This_stuffs_ �U  �M��U  �N��U  `O��U  �O��U  5#U/   �'U/      Appointment �� ��U  � ��U  Ы justforfun_justforfun_  ��U   � ��U  � ��U  �� ��U  `� ��U  �LU/   %KU/      Meeting     `���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �xU/   �xU/       Workout     Ѕ��U  ����U  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��U/   �U/       Some_stuffs ����U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �U/   )�U/      Meeting     `O��U  �O��U  �PSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  Pc��U  �U/   +�U/      Workout     �� ��U  @� ��U  �� justforfun_justforfun_  ��U  � ��U  Щ ��U  �� ��U  � ��U  qV/   IV/       Appointment �� ��U  P� ��U   � This_stuffs_This_stuffs_ �U  0� ��U  � ��U  �� ��U  p� ��U  L�`/   l�`/      Appointment                    justforfun_justforfun_                                       ��`/   ��`/       Birthday    �W��U  �X��U  `Yjustforfun_justforfun_ ��U  �[��U  `\��U   ]��U  �]��U  �a/   �a/       Meeting     �� ��U  P� ��U   � justforfun_justforfun_  ��U  0� ��U  � ��U  �� ��U  p� ��U  g7a/   �6a/       Meeting     P% ��U  & ��U  �) Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �8 ��U  `a/   �\a/       Meeting     `_ ��U   ` ��U  `d justforfun_justforfun_  ��U  �n ��U  Po ��U  �t ��U  �v ��U  ��a/   �a/      Workout     07��U  �7��U  p8justforfun_justforfun_ ��U  �:��U  0;��U  �;��U  p<��U  A�a/   �a/      Meeting     @� ��U   � ��U  �� justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U   ��U  ��a/   ��a/      Birthday    ����U  ���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �!b/   �"b/       Birthday    P#��U  $��U  �$justforfun_justforfun_ _ �U  �'��U   (��U  �(��U  �)��U  =rb/   kb/       Appointment ���U  ����U  оThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  W�b/   4�b/       Birthday    @��U  ���U  p�Some_stuffs_Some_stuffs_ �U  � ��U  ���U  0��U  ���U  #�b/   ��b/       Meeting     P���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  c/   �	c/       Meeting ent  ���U  ����U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  �/c/   =0c/      Birthday    P% ��U  & ��U  �) justforfun_justforfun_  ��U  P3 ��U  4 ��U  �7 ��U  �8 ��U  �[c/   �[c/      Appointment  � ��U  �� ��U  �� justforfun_justforfun_ _This_stuffs_This_stuffs_ �U   � ��U  �~c/   �~c/       Appointment  5��U  �5��U  �6This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `;��U  q�c/   ��c/       Meeting     �����U  p����U  p��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��c/   �c/       Appointment ����U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��c/   ��c/      Some_stuffs � ��U  � ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  & ��U  �d/   yd/       Workout     `���U  ����U  `�justforfun_justforfun_ ��U  ����U  `���U   ���U  ����U  
Ed/   7Fd/       Birthday    �� ��U  P� ��U   � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `� ��U  �gd/   �md/       Meeting ffs ����U  @���U  @This_stuffs_This_stuffs_ �U  p���U  0 ��U  � ��U  ���U  	�d/   ��d/      Birthday    P% ��U  & ��U  �) This_stuffs_This_stuffs_ �U  P3 ��U  4 ��U  �7 ��U  �8 ��U  8�d/   9�d/       Meeting     ����U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  ��d/   ��d/       Meeting     �s��U  Pt��U  �tThis_stuffs_This_stuffs_ �U  0w��U  �w��U  px��U  �x��U  �e/   te/      Meeting ent ���U  @��U   This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ��U  �)e/   %*e/      Birthday    0� ��U  � ��U  �� justforfun_justforfun_  ��U  P� ��U  � ��U  п ��U  �� ��U  �p/   ��o/      Workout �U  �+��U  p,��U  0-Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �1��U  �)p/   z%p/       Meeting      ��U  ���U  @�Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  @���U  =Pp/   �Pp/      Some_stuffs 0����U  �����U  P��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �����U  zp/   %zp/      Appointment �$��U  �%��U  P&Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   +��U  �p/   I�p/       Workout      ���U  ����U   �justforfun_justforfun_ ��U  `���U  ����U  ����U  `���U  x�p/   ��p/      Meeting     �� ��U  `� ��U   � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0� ��U  :�p/   T�p/      Some_stuffs P� ��U  p� ��U   � Some_stuffs_Some_stuffs_ �U   � ��U  � ��U  �� ��U  �� ��U  =q/   �q/       Birthday     ���U  ����U  @�justforfun_justforfun_ ��U  ����U  @���U   ���U  ����U  \=q/   L<q/       Meeting     0��U  ���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ��U  Jaq/   +_q/       Appointment �I��U  �J��U  `KSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �O��U  y�q/   j�q/       Birthday U  ���U  н��U  P�This_stuffs_This_stuffs_ �U  ���U  ����U  ����U  ���U  ��q/   ��q/      Meeting     �$��U  �%��U  P&This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   +��U  ��q/   4�q/       Birthday    �t��U  �u��U   vSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @z��U  Q�q/   	�q/       Some_stuffs p|��U  0}��U  �}This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Ё��U  
#r/   #r/       Birthday U  0���U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  �Kr/   3Hr/       Some_stuffs �� ��U  @� ��U  �� This_stuffs_This_stuffs_ �U  � ��U  Щ ��U  �� ��U  � ��U  sr/   rr/       Meeting      ���U  ����U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  ��r/   ��r/       Some_stuffs ����U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Џ��U  <�r/   C�r/      Some_stuffs 0���U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  5�r/   ��r/       Some_stuffs ���U  `���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  }s/   s/       Appointment �*��U  p+��U  0,Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �0��U  �6s/   87s/      Meeting �U  Ѕ��U  ����U  @�justforfun_justforfun_ ��U  `���U  ����U  `���U  ����U  P\s/   d\s/      Some_stuffs  ���U  ����U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0���U  t�s/   z�s/       Workout     p.��U  �.��U  p/Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  04��U  }�s/   l�s/       Meeting     ����U  @���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  t�s/   ~�s/      Appointment p� ��U  0� ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U   �s/   &�s/      Appointment ����U  P���U  �justforfun_justforfun_ _ �U  ����U  P���U  ���U  ����U  Lt/   & t/       Birthday    �t ��U  �v ��U  �z Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  �Kt/   �Lt/       Appointment @���U  ����U  @�This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  pt/   Znt/      Workout     @��U  ���U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  ��t/   �t/       Some_stuffs �� ��U  �� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   � ��U  �C/   BI/       Meeting     �Z ��U  p[ ��U  `_ Some_stuffs_Some_stuffs_ �U  pi ��U  0j ��U  �n ��U  Po ��U   g/   Dg/      Appointment P���U  ���U  лThis_stuffs_This_stuffs_ �U  P���U  ���U  ����U  ���U  3�/   ׏/       Workout ffs `���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  T�/   ^�/       Appointment ���U  ���U  P Some_stuffs_Some_stuffs_ �U  P#��U  $��U  �$��U  �%��U  R�/   ��/      Birthday U   ���U  ����U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  ��/   �/       Some_stuffs pi ��U  0j ��U  �n This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  �� ��U  {1�/   �2�/      Appointment `���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U   ���U  ����U  ����U  �U�/   �U�/      Some_stuffs �����U  @����U   ��justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  � ��U  @}�/   z}�/      Some_stuffs 0� ��U  � ��U  �� Some_stuffs_Some_stuffs_ �U  P� ��U  � ��U  п ��U  �� ��U  ���/   m��/       Appointment `O��U  �O��U  `PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �U��U  7ʀ/   �ƀ/       Appointment P ��U  !��U  �!Some_stuffs_Some_stuffs_ �U  �$��U  �%��U  P&��U  �1��U  ���/   ��/       Meeting ffs ���U  @��U  �This_stuffs_This_stuffs_ �U  P��U  ���U  ���U  ��U  H�/   ~�/      Workout      � ��U  �� ��U  @� This_stuffs_This_stuffs_ �U  �� ��U  P� ��U  � ��U  �� ��U  =�/   /A�/       Some_stuffs  o��U  �o��U   pThis_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  Pt��U  �g�/   h�/       Meeting     �T��U  0U��U  �Ujustforfun_justforfun_ _This_stuffs_This_stuffs_ �U  �Y��U  L��/   v��/      Appointment                    This_stuffs_This_stuffs_                                     ���/   流/       Workout ffs �����U  p����U  p��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ځ/   T��/       Appointment Pf��U  �f��U  Pgjustforfun_justforfun_ _ �U   i��U  �i��U   j��U  �j��U  \ �/   q �/       Birthday U  �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U  �'�/   �+�/       Some_stuffs `� ��U   � ��U  �� Some_stuffs_Some_stuffs_ �U  �� ��U  �� ��U  �� ��U  �� ��U  �O�/   �Q�/      Some_stuffs �
��U   ��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  �x�/   �x�/      Workout     �� ��U  P� ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p� ��U  �ɂ/   �Ƃ/       Appointment  ���U  ���U  `�Some_stuffs_Some_stuffs_ �U  ���U  ����U  ���U  ����U  ���/   ��/       Workout     ����U  `���U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  ��/   �/       Some_stuffs ���U   ��U  ��Some_stuffs_Some_stuffs_ �U   ���U  ����U  `���U   ���U  �>�/   �=�/       Some_stuffs ����U  `���U  ��justforfun_justforfun_ ��U  `���U  ����U  `���U  ����U  rc�/   1_�/       Some_stuffs 0� ��U  � ��U  �� Some_stuffs_Some_stuffs_ �U  �� ��U  P� ��U   � ��U  �� ��U  ���/   *��/       Birthday    �l��U  `m��U  �mSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �q��U  ��/   +��/       Workout     ����U  ���U  ��This_stuffs_This_stuffs_ �U  д��U  P���U  е��U  ����U  <؃/   _؃/      Meeting     ���U  `��U   Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ���U  ��/   ?��/       Workout     �����U  @����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  ^��/   ���/      Appointment �����U  @����U  ���Some_stuffs_Some_stuffs_ �U  �����U  P����U  �����U  @����U  �֎/   �Ў/      Meeting     `��U   ��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  �!�/   ��/       Meeting ffs ����U  `���U  ��This_stuffs_This_stuffs_ �U  `���U  ����U  ����U  `���U  �N�/   oJ�/       Birthday    ���U   ��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @��U  t�/   �m�/       Workout ent ����U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  ���/   ���/      Meeting     ����U  @���U   �This_stuffs_This_stuffs_ �U  ����U   ���U   ���U  ����U  ���/   쿏/       Meeting ent ���U  ����U  P�Some_stuffs_Some_stuffs_ �U  ����U  ���U  ����U  P���U  p�/   z�/       Meeting     �e��U  `f��U   gjustforfun_justforfun_ ��U  �i��U  `j��U   k��U  �k��U  ��/   ]�/      Workout     0��U  ���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  !��U  vW�/   AZ�/       Meeting     P���U  ����U  ��justforfun_justforfun_ _ �U  P���U  ���U  ����U  ����U  ���/   Æ�/       Workout     ���U  ����U  @�Some_stuffs_Some_stuffs_ �U  ����U   ���U  ����U  @���U  ��/   ��/       Meeting     0w��U  �w��U  pxSome_stuffs_Some_stuffs_ �U  pz��U  �z��U  p{��U  �{��U  l͐/   l͐/      Appointment @n��U  �n��U  @oThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @t��U  ,��/   0��/      Birthday nt ����U   ���U  ��justforfun_justforfun_ _ �U  ����U   ���U  ����U   ���U  ��/   !�/       Birthday nt е��U  ����U  �This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  @���U  pJ�/   	E�/      Meeting      ��U  ���U   Some_stuffs_Some_stuffs_ �U  ���U   ��U  ���U  @��U  �p�/   vp�/      Workout     � ��U  � ��U  � justforfun_justforfun_  ��U  0 ��U  � ��U  � ��U  � ��U  c��/   a��/       Workout      ��U  ���U  �justforfun_justforfun_ ��U   ��U  ���U  `��U  ���U  i��/   ���/      Some_stuffs ����U  P���U  �Some_stuffs_Some_stuffs_ �U  ����U  ����U  P���U  ����U  �	�/   ~�/       Workout     ����U  @���U  ��justforfun_justforfun_ ��U  @���U   ���U  ����U  ����U  �+�/   ,�/      Workout     �� ��U  P� ��U   � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p� ��U  �Z�/   Z�/       Workout     p.��U  �.��U  p/justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  04��U  �~�/   \~�/      Workout �U  �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U  ���/   ϥ�/      Some_stuffs ����U  @���U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  RΒ/   /ϒ/       Meeting     �	��U  �
��U  `justforfun_justforfun_ ��U   ��U  ���U  ���U  `��U  `��/   ���/       Meeting     ���U  ���U  `Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U   
��U  �ĝ/   ŝ/      Appointment  ���U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  ��/   ��/      Appointment �� ��U  `� ��U   � This_stuffs_This_stuffs_ �U  0� ��U  � ��U  p� ��U  0� ��U  ��/   ��/       Meeting      x��U  �x��U  �yjustforfun_justforfun_ ��U   |��U  �|��U  �}��U  @~��U  �d�/   dh�/       Appointment `���U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  ���/   b��/       Birthday    ����U  ����U   �Some_stuffs_Some_stuffs_ �U  ����U   ���U  ����U  ����U  0��/   g��/      Workout     �����U  `����U  ��justforfun_justforfun_ ���U  �����U  p����U  0����U  ����U  ���/   ��/       Birthday    @���U  ����U  @�This_stuffs_This_stuffs_ �U  @���U  ����U  @���U  ����U  �)�/   l*�/      Some_stuffs  � ��U  �� ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   � ��U  �u�/   �z�/       Some_stuffs ���U  `��U   justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ���U  Ԝ�/   �/      Meeting     Б��U  P���U  ВSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  ş/   �ɟ/       Workout     �E��U  `F��U   GThis_stuffs_This_stuffs_ �U  �U��U  pV��U  �I��U  �J��U  ��/   
�/      Appointment ���U  ���U  P This_stuffs_This_stuffs_ �U  P#��U  $��U  �$��U  �%��U  ��/   ��/       Some_stuffs �+��U  �,��U   -This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �0��U  5<�/   �=�/      Birthday    �]��U  p^��U  0_Some_stuffs_Some_stuffs_ �U  0b��U  �b��U  �c��U  Pd��U  �`�/   ya�/       Some_stuffs �;��U  p<��U  �<Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p@��U  ���/   ͌�/      Workout     0����U  ����U  ���This_stuffs_This_stuffs_ �U   ����U  �����U  �����U  p����U  㭠/   ��/       Meeting     P���U  ���U  БThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  q��/   L��/      Some_stuffs @���U   ���U  ��Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ���U  �(�/   )�/       Birthday    �� ��U   ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  �q�/   �p�/       Workout     �y��U  @z��U  �zThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  |��/   ���/      Meeting     �:��U  0;��U  �;justforfun_justforfun_ ��U  �=��U  p>��U  �>��U  p?��U  ��/   ��/      Some_stuffs ����U  ����U  P�Some_stuffs_Some_stuffs_ �U  ����U  @���U   ���U  ����U  09�/   79�/      Birthday    `���U   ���U  ��This_stuffs_This_stuffs_ �U  `���U  ����U  ����U   ���U   Z�/   :Z�/      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��/   �	�/      Some_stuffs  5��U  �5��U   6This_stuffs_This_stuffs_ �U  �8��U  @9��U  `R��U   S��U  E.�/   I4�/       Appointment  =��U  �=��U  `2justforfun_justforfun_ ��U   5��U  �5��U  �6��U   7��U  ��/   ���/      Some_stuffs ���U  p��U  0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ~��/   詭/       Some_stuffs  ���U  ����U  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  F��/   ��/       Birthday     ��U  ���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ��U  ��/   M�/       Some_stuffs P����U  ����U  P��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  -E�/   �F�/       Birthday    p���U  0���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  �g�/   ]o�/      Birthday    ����U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ��/   I��/      Meeting                        Some_stuffs_Some_stuffs_                                     ���/   M��/       Workout  U  �
��U   ��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @��U  �߮/    �/       Appointment �Z��U   [��U  �[justforfun_justforfun_ ��U  �^��U   _��U  �_��U  �`��U  ��/   ��/      Meeting �U  p\��U  0]��U  �]Some_stuffs_Some_stuffs_ �U  �`��U  pa��U  0b��U  �b��U  �-�/   �.�/      Workout     P% ��U  & ��U  �) justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  �8 ��U  U�/   �V�/      Some_stuffs ����U  @���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  i��/   /      Workout     `!��U  �!��U   :Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �&��U  	��/   ��/       Appointment �� ��U  @� ��U   � justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  P� ��U  }�/   :�/      Birthday fs �L��U  `M��U  �MSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �l��U  5@�/   A�/      Appointment 0� ��U  � ��U  p� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0� ��U   j�/   j�/       Some_stuffs ���U  ����U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ���/   D��/       Meeting     �l��U  Pm��U  �mThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �q��U  ׳�/   ���/       Some_stuffs �S ��U  �U ��U  �Z justforfun_justforfun_  ��U  `d ��U   e ��U  pi ��U  0j ��U  I۰/   �ް/      Birthday    ���U  `���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  #�/   ���/       Appointment �2��U  @3��U  �3Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U   8��U  )�/   (�/      Meeting      ��U  ���U  �BThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  �#��U  �u�/   �z�/       Meeting �U  0���U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �Q�/   �K�/       Workout     �F��U  0G��U  �GThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �K��U  �p�/   Tq�/       Birthday    л��U  ����U  �Some_stuffs_Some_stuffs_ �U  ����U  ���U  ���U  ����U  5��/   b��/      Birthday    ����U  @���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  ��/   �/       Workout     �����U  p����U  p��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  \�/   ��/      Some_stuffs �� ��U  p� ��U  0� This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  �� ��U  A;�/   �9�/       Birthday    p� ��U  0� ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  0_�/   X_�/       Birthday    `� ��U   � ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  ���/   1��/      Birthday    �V��U  �W��U  pXjustforfun_justforfun_ ��U  0[��U  �[��U  p\��U  0]��U  ��/   `��/       Birthday    ����U   ���U  p�justforfun_justforfun_ ��U  p���U  ���U  ����U  @���U  �ӽ/   �׽/      Some_stuffs `���U   ���U  ��justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  ����U  ��/   ���/       Workout ffs `���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  I#�/   �"�/      Appointment ����U  @���U   �justforfun_justforfun_ ��U  ����U  0���U  ����U  p���U  �I�/   �J�/       Birthday    �� ��U  �� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   � ��U  hq�/   �q�/       Appointment �B��U  `C��U   DSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �H��U  њ�/   +��/       Some_stuffs `���U  ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  R��/   ���/       Appointment �s��U  @t��U  �tThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �x��U  ��/   B�/       Appointment ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  ����U  `���U   ���U  U�/   
�/       Workout     ���U  ����U  @�Some_stuffs_Some_stuffs_ �U  @���U  ����U  @���U  ����U  7�/   G5�/       Appointment  ��U  ���U  `justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U   ��U  EX�/   �[�/       Birthday    �'��U   (��U  �(This_stuffs_This_stuffs_ �U  �+��U  �,��U   -��U  �-��U  ؂�/   邿/      Workout     `Y��U  �Y��U  �Zjustforfun_justforfun_ ��U   ]��U  �]��U  �^��U   _��U  �п/   �ο/      Appointment @���U   ���U  ��This_stuffs_This_stuffs_ �U  @���U  ����U  ����U   ���U  L��/   ���/      Workout      ��U  ���U  @Some_stuffs_Some_stuffs_ �U  @��U   ��U  ���U  ���U  ��/   ��/      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             nC�/   �I�/      Meeting     �a��U  Pb��U  �bThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �f��U  l�/   �j�/       Workout      ��U  ���U  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  e��/   ��/       Birthday    ���U  Џ��U  P�Some_stuffs_Some_stuffs_ �U  В��U  ����U  ���U  ����U  ���/   ���/       Birthday    p���U  0���U  ��This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  P���U  �T
 /   �U
 /       Appointment �@ ��U  �A ��U  pE This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  �U ��U  ?~
 /   '}
 /       Appointment 0_��U  �_��U  �`Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �e��U  ߦ
 /   l�
 /       Some_stuffs 0a��U  �a��U  0bSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   g��U  �
 /   <�
 /      Some_stuffs � ��U  � ��U  � justforfun_justforfun_  ��U  0 ��U  � ��U  � ��U  � ��U  ��
 /   �
 /       Appointment P����U  ����U  P��This_stuffs_This_stuffs_ �U  P����U  ����U  �����U  @����U  ' /   j /       Workout �U  �>��U  p?��U  �?Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  �D��U  �B /   �B /       Appointment ����U  ���U  ��justforfun_justforfun_ ��U  е��U  ����U  ���U  ����U  $c /   Oc /      Meeting     �����U  `����U  ��Some_stuffs_Some_stuffs_ �U  �����U  p����U  0����U  ����U  � /   � /       Some_stuffs Ю��U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  � /   � /      Some_stuffs 0� ��U  � ��U  �� Some_stuffs_Some_stuffs_ �U  �� ��U  P� ��U   � ��U  �� ��U  �� /   �� /       Appointment �� ��U  �� ��U  @� justforfun_justforfun_ ��U  �� ��U  @ ��U   ��U  ���U  �  /   � /       Some_stuffs ����U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  0) /   k) /      Meeting �U  �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U  �S /   �M /      Meeting     `K��U   L��U  �LSome_stuffs_Some_stuffs_ �U  `O��U  �O��U  �P��U  `Q��U  �v /   �u /      Workout     м ��U  �� ��U  P� This_stuffs_This_stuffs_ �U  P� ��U  � ��U  �� ��U  �� ��U  ٣ /   �� /       Appointment  ��U  ���U   justforfun_justforfun_ ��U  ���U   ��U  ���U  @��U  �� /   �� /      Birthday    �����U  p����U  p��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �� /   9� /      Meeting ent P% ��U  & ��U  �) justforfun_justforfun_ _ �U  P3 ��U  4 ��U  �7 ��U  �8 ��U  	 /   ^ /       Some_stuffs Ю��U  P���U  �Some_stuffs_Some_stuffs_ �U  ���U  ����U  `���U   ���U  w9 /   �> /       Some_stuffs �$��U  �%��U  P&This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   +��U  4e /   :e /       Meeting     �Z ��U  p[ ��U  `_ justforfun_justforfun_  ��U  pi ��U  0j ��U  �n ��U  Po ��U  �� /   s� /       Meeting     �_��U  �`��U   aSome_stuffs_Some_stuffs_ �U  �c��U  `d��U  �d��U  `e��U  �� /   I� /       Workout     @���U   ���U  ��Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ����U  �� /   �� /       Birthday    �� ��U  �� ��U   � justforfun_justforfun_  ��U  p� ��U  �� ��U   � ��U  �� ��U  6� /   �� /       Appointment 0���U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `���U  �* /   �* /       Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �Q /   �J /       Some_stuffs �����U  p����U  p��This_stuffs_This_stuffs_ �U  @����U  ����U  P����U  ����U  p /   �r /      Meeting     @���U  ����U  @�This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U   ���U  � /   Ě /       Meeting ffs  ���U  ����U  `�justforfun_justforfun_ ��U  ����U  `���U   ���U  ����U  P� /   v� /      Some_stuffs @���U   ���U  ��This_stuffs_This_stuffs_ �U  @���U  ����U  ����U  @���U  � /   A� /       Some_stuffs @7��U   8��U  �8Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   =��U  P� /   �� /      Workout �U  @� ��U   � ��U  �� justforfun_justforfun_  ��U  � ��U  �� ��U  �� ��U  P� ��U  �� /   �� /       Some_stuffs �`��U  pa��U  0bSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �f��U  X /   s /      Appointment @��U   ��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �
��U  h8 /   }8 /      Birthday U  �����U  �����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @����U  �V /   e\ /       Appointment �E��U  `F��U   GSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �J��U  �~ /   [� /       Appointment ���U  p���U  �This_stuffs_This_stuffs_ �U  0���U  ���U  ����U  p���U  �� /   � /       Appointment @� ��U   � ��U  �� This_stuffs_This_stuffs_ �U   ��U  ���U  @��U   ��U  �� /   �� /       Meeting �U  �W��U  pX��U  �Xjustforfun_justforfun_ ��U  0[��U  �[��U  0\��U  �\��U  X� /   �� /       Workout �U  �����U  �����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @����U  ~ /   � /       Workout ent @��U  ���U  `Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  @��U  �G /   (D /       Workout ffs @���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  �o /   Pq /       Some_stuffs �l��U  Pm��U  �mSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �q��U  � /   �� /      Appointment �t��U  �u��U   vSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �z��U  e� /   �� /       Birthday    ���U  ����U  �justforfun_justforfun_ ��U  г��U  ����U  ���U  ����U  �� /   ,� /       Some_stuffs �� ��U  P� ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p� ��U  � /   F /       Appointment ����U  ����U  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �+ /   �3 /       Birthday    ���U  ���U  @Some_stuffs_Some_stuffs_ �U  ���U  0��U  ���U  `	��U  (X /   [X /       Some_stuffs `{��U  �{��U  �|justforfun_justforfun_ ��U  ���U   ���U  ����U  `���U  ~| /   r� /      Birthday    `O��U  �O��U  �PSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  Pc��U  �� /   �� /      Appointment  J ��U  �J ��U  �N This_stuffs_This_stuffs_ �U  �Z ��U  p[ ��U  `_ ��U   ` ��U  � /   +� /       Some_stuffs ���U  ���U    This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p$��U  � /   �� /       Birthday nt �<��U  p=��U  �=This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �A��U   /   " /      Meeting     �O��U  pP��U  �PSome_stuffs_Some_stuffs_ �U  pS��U  0T��U  �T��U  0U��U  ? /   IB /       Meeting �U  ����U  P���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  Le /   Qe /      Some_stuffs ���U  ���U  pSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  p��U  '� /   � /       Meeting      ��U  ���U  �	Some_stuffs_Some_stuffs_ �U  �"��U  @#��U  ���U  `��U  � /   #� /      Workout     ����U  ����U  �justforfun_justforfun_ _ �U  ����U  ����U   ���U  ����U  >�( /   n�( /       Birthday    ����U  ����U  @�This_stuffs_This_stuffs_ �U  ����U   ���U  п��U  P���U  )) /   @%) /      Workout     D��U  �D��U  PESome_stuffs_Some_stuffs_ �U  �G��U  �H��U   I��U  �I��U  �S) /   T) /       Birthday U  ���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �t) /   �r) /      Meeting     P����U  ����U  P��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @����U  ҝ) /   ��) /       Some_stuffs �����U  �����U  ���justforfun_justforfun_ _ his_stuffs_This_stuffs_ �U  @����U  ��) /   h�) /       Birthday    @��U   ��U  �This_stuffs_This_stuffs_ �U  ���U  ���U   ��U  ���U  M* /   ~* /       Appointment ����U  p���U  ��This_stuffs_This_stuffs_ �U  ����U  ����U  0���U  ����U  �6* /   `;* /       Meeting      6��U  �6��U  @7This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �;��U  Ad* /   d* /       Some_stuffs  ���U  ����U    justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ���U  ^�* /   p�* /       Appointment `Y��U  �Y��U  �ZSome_stuffs_Some_stuffs_ �U   ]��U  �]��U  �^��U   _��U  ��* /   ��* /      Workout     ���U  `���U   �This_stuffs_This_stuffs_ �U  ���U  `���U   ���U  ���U  Q�* /   <�* /       Meeting     `>��U  �>��U  �?This_stuffs_This_stuffs_ �U  �B��U  `C��U   D��U  �D��U  �+ /   ��* /       Workout     P���U  ���U  лSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  $+ /   � + /       Some_stuffs o��U  �o��U  �~justforfun_justforfun_ ��U  `r��U   s��U  �s��U  `t��U  TJ+ /   �J+ /      Appointment `� ��U   � ��U  �� Some_stuffs_Some_stuffs_ �U  �� ��U  `� ��U  p� ��U  �� ��U  �m+ /    n+ /      Meeting     ����U  ����U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  ��+ /   Q�+ /       Some_stuffs P% ��U  & ��U  �) Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �8 ��U  5�+ /   0�+ /       Workout     �� ��U  p� ��U  0� justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  @� ��U  E�+ /   ��+ /      Birthday    ����U  ����U   �This_stuffs_This_stuffs_ �U  ����U  `���U   ���U  ����U  !
, /   �, /       Workout     p���U  0���U  ��This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  0���U  7, /   �1, /       Meeting     ����U   ���U  ��This_stuffs_This_stuffs_ �U  ����U   ���U  ����U   ���U  �X, /   �`, /       Appointment `K��U   L��U  �LSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `Q��U  �, /   )�, /      Birthday    �(��U  p)��U  �)This_stuffs_This_stuffs_ �U  0,��U  �,��U  p-��U  0.��U  ��, /   ��, /       Birthday    ���U  ���U    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p$��U  e�, /   ��, /       Some_stuffs �� ��U  �� ��U  0� This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  � ��U  � - /   � - /      Meeting     ���U  ���U    Some_stuffs_Some_stuffs_ �U   :��U  �:��U  �#��U  p$��U  �B- /   E- /      Appointment ���U  ����U  оThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  `n- /   }n- /      Birthday    `w��U  �w��U  �xjustforfun_justforfun_ ��U  `{��U  �{��U  �|��U  `}��U  8 /   8 /       Birthday    ����U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  �?8 /   �?8 /      Meeting     @���U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  �j8 /   k8 /       Meeting     �� ��U  � ��U  Ы This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `� ��U  c�8 /   ��8 /       Some_stuffs  ;��U  �;��U  �<justforfun_justforfun_ ��U  `?��U  �?��U  `@��U   A��U  f�8 /   o�8 /       Meeting     �� ��U  �� ��U  P� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   � ��U  ��8 /   ��8 /       Meeting ffs �����U  p����U  p��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �,9 /   #29 /       Some_stuffs �� ��U  @� ��U  �� justforfun_justforfun_  ��U  � ��U  Щ ��U  �� ��U  � ��U  !R9 /   �W9 /      Meeting �U   � ��U  �� ��U  �� This_stuffs_This_stuffs_ �U   � ��U  �� ��U  @� ��U   � ��U  }}9 /   z9 /      Birthday    �_��U  �`��U   aSome_stuffs_Some_stuffs_ �U  �c��U  `d��U  �d��U  `e��U  С9 /   ��9 /      Some_stuffs �t ��U  �v ��U  �z This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  <�9 /   W�9 /       Workout     ���U  `���U   �Some_stuffs_Some_stuffs_ �U  ����U  `���U  ���U  ����U  �: /   �: /       Meeting     �� ��U  P� ��U   � Some_stuffs_Some_stuffs_ �U  0� ��U  � ��U  �� ��U  p� ��U  =?: /   eA: /       Birthday    �� ��U  � ��U  Ы This_stuffs_This_stuffs_ �U   � ��U  � ��U  �� ��U  `� ��U  �c: /   �g: /       Workout     p� ��U  0� ��U  �� Some_stuffs_Some_stuffs_ �U  �� ��U  0� ��U  м ��U  �� ��U  h�: /   h�: /       Workout     ����U  @���U  ��Some_stuffs_Some_stuffs_ �U  ����U  @���U   ���U  ����U  ��: /   ı: /      Birthday    �:��U  `;��U   <This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �A��U  p�: /   r�: /       Appointment ���U  ����U  P�Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ����U  I; /   ��: /      Workout     P��U   ��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `��U  f*; /   u%; /       Workout     `2��U   3��U  �3This_stuffs_This_stuffs_ �U  �6��U   7��U  �7��U  �8��U  1T; /   �S; /      Meeting     �X��U   Y��U  �YThis_stuffs_This_stuffs_ �U  �[��U  0\��U  �\��U  0]��U  gu; /   cy; /       Meeting ent  ��U  ���U  �justforfun_justforfun_ _ �U   ��U  ���U  `��U  ���U  2�; /   ��; /       Birthday    p+��U  �+��U  p,This_stuffs_This_stuffs_ �U  �.��U  p/��U  �/��U  p0��U  ��; /   ��; /       Appointment �:��U  `;��U   <This_stuffs_This_stuffs_ �U  �?��U  `@��U   A��U  �A��U  ��; /   %�; /       Birthday U  0<��U  �<��U  p=This_stuffs_This_stuffs_ �U  �?��U  0@��U  �@��U  `A��U  a< /   �< /       Workout ffs � ��U  Щ ��U  �� This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  � ��U  ,�< /   P�< /      Appointment �����U  @����U  ���This_stuffs_This_stuffs_ �U  �����U  P����U  �����U  @����U  ~[G /   �`G /      Meeting      � ��U  �� ��U  @� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  k�G /   �G /       Birthday    p���U  ���U  ��This_stuffs_This_stuffs_ �U  ���U  ����U  ���U  ����U  L�G /   ~�G /       Birthday    �
��U   ��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ��U  ��G /   ��G /      Appointment p���U  0���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0���U  	�G /   ��G /       Workout     ����U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  iH /   �!H /       Meeting     � ��U  ���U  0Some_stuffs_Some_stuffs_ �U  ���U  ���U   ��U  ���U  �JH /   IH /       Some_stuffs �F��U  �G��U  `Hjustforfun_justforfun_ ��U  `K��U   L��U  �L��U  `M��U   rH /   rH /       Appointment �(��U  P)��U  �)This_stuffs_This_stuffs_ �U  �+��U  p,��U  0-��U  �-��U  ��H /   O�H /       Workout     ����U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U  ����U   ���U  ����U  0�H /   )�H /       Workout     ����U  ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��H /   D�H /       Birthday    �t��U  �u��U   vThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @z��U  [
I /   �
I /       Meeting     ����U  p���U  ��Some_stuffs_Some_stuffs_ �U  @���U   ���U  ����U   ���U  �4I /   �4I /      Workout      v��U  �v��U  `wThis_stuffs_This_stuffs_ �U  �y��U  �z��U  `{��U  �{��U  MWI /   �WI /      Meeting     �� ��U  �� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `� ��U  t�I /   1~I /       Appointment ����U  ����U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  
�I /   A�I /      Workout     �*��U  p+��U  0,Some_stuffs_Some_stuffs_ �U  �.��U  p/��U  �/��U  �0��U  :�I /   Y�I /       Some_stuffs  0��U  �0��U   =This_stuffs_This_stuffs_ �U  �3��U  �4��U   5��U  �5��U  �I /   =�I /      Birthday    � ��U  � ��U  � justforfun_justforfun_  ��U   ! ��U  �! ��U  P% ��U  & ��U  �J /   �J /      Appointment ����U  `���U   �Some_stuffs_Some_stuffs_ �U  ����U  `���U  ����U  `���U  �EJ /   �@J /       Appointment ����U  @���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �gJ /   �oJ /       Workout     �� ��U  @ ��U   Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  ��J /   =�J /       Meeting     p��U  ���U  �Some_stuffs_Some_stuffs_ �U  ���U   '��U  P��U  ��U  (�J /   <�J /      Appointment �� ��U  �� ��U  P� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   � ��U   �J /   �J /      Appointment p� ��U  �� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   � ��U  �K /   $K /       Some_stuffs p\��U  0]��U  �]Some_stuffs_Some_stuffs_ �U  �`��U  pa��U  0b��U  �b��U  �-K /   �1K /       Appointment ����U  P���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  �SK /   �SK /       Appointment ����U   ���U  ��Some_stuffs_Some_stuffs_ �U  `���U   ���U  ����U  ����U  �K /   C�K /       Workout     �~��U   ��U  �pSome_stuffs_Some_stuffs_ �U  �s��U  `t��U  �t��U  �u��U  ��K /   ��K /       Meeting ent p9��U  0:��U  �:Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p>��U  ��K /   x�K /       Workout     �� ��U  �� ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  P�K /   _�K /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             a�V /   ��V /       Workout     ����U  ����U  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��V /   /�V /       Some_stuffs  w��U  �w��U   xSome_stuffs_Some_stuffs_ �U  �z��U  �{��U   |��U  �|��U  ��V /   ��V /       Birthday nt �m��U  Pn��U  oSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   s��U  �9W /   J=W /       Appointment �����U  @����U  ���This_stuffs_This_stuffs_ �U  �����U  P����U  �����U  @����U  xhW /   xhW /       Workout     `� ��U   � ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  ͌W /   ^�W /      Workout     ����U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��W /   S�W /       Appointment �k��U  l��U  �ljustforfun_justforfun_ ��U  o��U  �o��U  �~��U   ��U  ��W /   Z�W /      Birthday    ����U  0���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  � X /   �W /       Birthday    ����U  P���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  cMX /   �LX /       Workout     ����U  ���U  гjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  P���U   vX /   5vX /       Workout     j��U  �j��U  �kThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �o��U  �X /   Y�X /      Appointment  H��U  �H��U  �UThis_stuffs_This_stuffs_ �U  `K��U   L��U  �L��U  `M��U  ��X /   ��X /       Some_stuffs 0[��U  �[��U  p\This_stuffs_This_stuffs_ �U  0_��U  �_��U  �`��U  pa��U  ��X /    �X /       Workout     p���U  0���U  ��This_stuffs_This_stuffs_ �U  ����U  ����U  p���U  P���U  yY /   LY /       Workout     Pf��U  �f��U  Pgjustforfun_justforfun_ ��U   i��U  �i��U   j��U  �j��U  �<Y /   �7Y /       Appointment � ��U  � ��U  � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  � ��U  TbY /   ebY /      Meeting �U  `r��U   s��U  �sSome_stuffs_Some_stuffs_ �U   v��U  �v��U  `w��U  �w��U  �Y /   ��Y /      Birthday    � ��U  Щ ��U  �� Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  � ��U  ҩY /   �Y /       Appointment �I��U  �J��U  `KThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �O��U  �Y /   2�Y /      Appointment �� ��U  @� ��U  �� This_stuffs_This_stuffs_ �U  � ��U  Щ ��U  �� ��U  � ��U  ��Y /   ��Y /       Some_stuffs p6��U  07��U  �7This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �;��U  �"Z /   �"Z /      Birthday    �'��U  p(��U  �(This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �,��U  @GZ /   %KZ /      Birthday fs �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U  vZ /   LmZ /       Birthday    д��U  P���U  еSome_stuffs_Some_stuffs_ �U  P���U   ���U  ����U  @���U  �Z /   ��Z /      Workout     �3��U  p4��U  �4Some_stuffs_Some_stuffs_ �U  �7��U  08��U  �8��U  p9��U  =�Z /   /�Z /       Workout     �*��U  p+��U  0,Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �0��U  ��Z /   ��Z /       Workout     0����U  ����U  ���Some_stuffs_Some_stuffs_ �U   ����U  �����U  �����U  p����U  �[ /   ?[ /       Workout      R��U  �R��U  `SThis_stuffs_This_stuffs_ �U  �V��U  �W��U  pX��U  0Y��U  ��e /   ��e /      Appointment ����U  ����U  `�justforfun_justforfun_ ��U  `���U  ����U  ����U   ���U  �f /   �f /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �5f /   �5f /       Some_stuffs �h��U  �i��U  jThis_stuffs_This_stuffs_ �U  �l��U  Pm��U  �m��U  Pn��U  eTf /   �Yf /       Workout     �� ��U  @ ��U   Some_stuffs_Some_stuffs_ �U  ���U  ���U  @��U   ��U  u{f /   3}f /      Meeting ffs ���U  @��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ��U  ��f /   ȣf /      Appointment  J ��U  �J ��U  �N justforfun_justforfun_  ��U  �Z ��U  p[ ��U  `_ ��U   ` ��U  P�f /   \�f /       Workout �U   0��U  �0��U   =This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �5��U  ��f /   ��f /       Birthday nt @���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  �g /   wg /      Appointment   ��U  � ��U   ! Some_stuffs_Some_stuffs_ �U  �) ��U  P* ��U  �. ��U  �/ ��U  �?g /   @g /       Some_stuffs �A��U  �B��U   Cjustforfun_justforfun_ ��U  �E��U  `F��U  �F��U  �G��U  .hg /   0gg /       Meeting     �z��U   {��U  �{This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P��U  ^�g /   Ւg /      Appointment ���U  @��U  �This_stuffs_This_stuffs_ �U   ��U  ���U   ��U  ���U  ��g /   ��g /      Appointment  � ��U  �� ��U  �� This_stuffs_This_stuffs_ �U  �� ��U  p� ��U  �� ��U  P� ��U  )h /   �	h /      Meeting �U  �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U  /h /   �)h /       Some_stuffs ���U   ��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  6Ph /   7Th /      Workout ent ����U  P���U  ��This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  Fwh /   Zyh /       Appointment  ���U  ����U  @�Some_stuffs_Some_stuffs_ �U  ����U  ����U  @���U   ���U  ¥h /   �h /       Meeting     �� ��U  �� ��U  P� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   � ��U  >�h /   s�h /       Birthday    �W��U  pX��U   YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �]��U  �i /   yi /       Appointment P���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  Bi /   `?i /       Workout     ����U  ���U  ��This_stuffs_This_stuffs_ �U  ����U  P���U  ����U  ����U  gi /   �gi /       Workout     p���U  0���U  ��This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ���U  ��i /   "�i /       Birthday nt p���U  ����U  p�justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  `���U  h�i /   j�i /      Some_stuffs p\��U  0]��U  �]Some_stuffs_Some_stuffs_ �U  �`��U  pa��U  0b��U  �b��U  B�i /   D�i /       Appointment D��U  �D��U  PEjustforfun_justforfun_ ��U  �G��U  �H��U   I��U  �I��U  ij /   A�i /      Workout      v��U  �v��U  `wSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �{��U  �$j /   �$j /      Workout ffs ����U  P���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  %Oj /   ~Nj /       Birthday nt �� ��U  @� ��U  `� This_stuffs_This_stuffs_ �U   � ��U  �� ��U  �� ��U  `� ��U  �yj /   �wj /       Some_stuffs ���U  `��U  �Some_stuffs_Some_stuffs_ �U  ���U  ���U    ��U  � ��U  �"u /   �"u /      Birthday     0��U  �0��U   =Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �5��U  �Ku /   �Lu /       Appointment Ё��U  p���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �ou /   �tu /       Workout     p���U  ����U  p�Some_stuffs_Some_stuffs_ �U  0��U  ���U  ���U  `��U  5�u /   �u /       Workout     �t ��U  �v ��U  �z This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  ��u /   �u /      Some_stuffs �� ��U  @� ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  � ��U  �u /   :�u /      Birthday     A��U  �A��U  �Bjustforfun_justforfun_ ��U  �E��U  `F��U   G��U  �G��U   v /   v /       Appointment ���U  `��U   This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  �5v /   �7v /      Appointment e��U  �e��U  fThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �j��U  	_v /   �[v /      Birthday U  p���U  P���U  �Some_stuffs_Some_stuffs_ �U  Б��U  P���U  В��U  ����U  �v /   �v /      Appointment ���U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  ��v /   �v /      Workout     ����U  ����U  �Some_stuffs_Some_stuffs_ �U  ����U  P���U  ���U  ����U  d�v /   ��v /       Workout     02��U  �2��U  �3Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �7��U  �v /   1�v /      Some_stuffs `U��U  �U��U  �VThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   [��U  w /   �w /       Some_stuffs ����U  ����U  p�This_stuffs_This_stuffs_ �U  P���U  ���U  Б��U  P���U  �Jw /   lDw /       Workout     �� ��U  � ��U  Ы This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `� ��U  �nw /   �nw /      Some_stuffs                    justforfun_justforfun_                                       �w /   x�w /       Workout     ����U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  A�w /   '�w /       Birthday    �Y��U  �Z��U  0[This_stuffs_This_stuffs_ �U  �]��U  p^��U  0_��U  �_��U  $�w /   )�w /       Meeting  nt  ���U  ����U   �Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ����U  �x /   0x /       Meeting     `���U  ���U  ��justforfun_justforfun_ _ his_stuffs_This_stuffs_ �U  б��U  F0x /   �3x /       Birthday    �
��U   ��U  �justforfun_justforfun_ ��U   ��U  ���U  @��U   ��U  ]^x /   �\x /      Appointment ���U  p���U  �justforfun_justforfun_ _ �U  0���U  ���U  ����U  p���U  q|x /   �|x /       Meeting      ��U  ���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pC��U  ��x /   ޥx /       Appointment   ��U  � ��U  `!This_stuffs_This_stuffs_ �U  �#��U  p$��U  0%��U  �%��U  (�x /   Y�x /       Some_stuffs p� ��U  0� ��U  �� This_stuffs_This_stuffs_ �U  �� ��U  0� ��U  м ��U  �� ��U  ��x /   ��x /      Birthday fs P���U  У��U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �y /   � y /       Appointment p���U  0���U  ��justforfun_justforfun_ ��U  ����U  ����U  p���U  P���U  �@y /   �@y /       Birthday    `K��U   L��U  �LSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `Q��U  6gy /   hoy /       Workout     0 ��U  � ��U  � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �! ��U  �y /   N�y /       Appointment 06��U  �6��U  07This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0;��U  �y /   Ļy /       Some_stuffs ���U  И��U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  �d� /   �j� /      Some_stuffs �H��U  PI��U  JSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �M��U  ��� /   ��� /       Birthday    `���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��� /   ʷ� /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �ۄ /   #�� /       Meeting     �t��U  �u��U   vjustforfun_justforfun_ ��U  �x��U  `y��U  �y��U  �z��U  (� /   b� /      Meeting �U  Pg��U  h��U  �hThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Pm��U  0(� /   b(� /      Meeting     @���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  �S� /   �S� /      Some_stuffs �y��U  �z��U  `{justforfun_justforfun_ ��U  ����U  p���U  ���U   ���U  �z� /   y� /       Appointment �� ��U  P� ��U  � justforfun_justforfun_  ��U  0� ��U  �� ��U  �� ��U  p� ��U  u�� /   %�� /       Birthday    P���U  ���U  Бjustforfun_justforfun_ ��U  ���U  ����U  P���U  ���U  eƅ /   ZɅ /       Appointment �� ��U  P� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p� ��U  � /   ,� /      Workout     Pf��U  �f��U  Pgjustforfun_justforfun_ ��U   i��U  �i��U   j��U  �j��U  z� /   �� /      Birthday    ����U  @���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  5;� /   �:� /       Meeting      ���U  ����U   �Some_stuffs_Some_stuffs_ �U  @���U   ���U  ����U  @���U  Bb� /   �`� /       Some_stuffs p|��U  0}��U  �}This_stuffs_This_stuffs_ �U  P���U  Ѐ��U  P���U  Ё��U  8�� /   C�� /       Meeting     л��U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  5�� /   ��� /       Meeting     ����U  `���U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �׆ /   :Ն /       Workout     ����U  @���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  z)� /   �'� /       Workout �U  ����U  @���U  ��justforfun_justforfun_ ��U  @���U   ���U  ����U  0���U  �P� /   {K� /       Workout     @��U  ���U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  �r� /   q� /      Workout     `!��U  �!��U   :justforfun_justforfun_ ��U  0%��U  �%��U  p&��U  �&��U  �� /   ș� /       Some_stuffs  ���U  ����U  P�Some_stuffs_Some_stuffs_ �U  ����U   ���U  ����U  0���U  @�� /   y�� /      Birthday     � ��U  �� ��U  �� justforfun_justforfun_  ��U   � ��U  �� ��U  @� ��U   � ��U  D� /   g� /      Meeting     ����U  p���U  �Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   ���U  W� /   G� /       Birthday    p���U  0���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �8� /   �8� /       Birthday    @� ��U   � ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  �^� /   �[� /       Workout �U  P���U  ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  П��U  �� /   H�� /      Meeting     ���U  ���U    This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p$��U  Ы� /   k�� /       Meeting     P� ��U  @� ��U  0� justforfun_justforfun_  ��U  0� ��U  �� ��U  �� ��U  p� ��U  �؈ /   �؈ /      Meeting                        This_stuffs_This_stuffs_                                     �� /   �� /      Appointment �����U  @����U   ��justforfun_justforfun_ ���U  �����U  �  ��U  � ��U  � ��U  �Г /   &ԓ /       Appointment ���U  ����U  ��justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ���U  J�� /   o�� /       Workout     ����U   ���U  p�Some_stuffs_Some_stuffs_ �U  p���U  ���U  ����U  @���U  Q� /   :!� /       Appointment  <��U  �<��U  `>Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `C��U  �j� /   �j� /       Some_stuffs ����U  @���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �� /   )�� /       Birthday    ����U  p���U  0�justforfun_justforfun_ ��U  ����U  p���U  ����U  ����U  ��� /   ��� /       Some_stuffs  ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  �� /   �� /      Some_stuffs P����U  ����U  @��justforfun_justforfun_ _ �U  P����U  �����U  0����U  �����U  b� /   I� /       Meeting     ����U  ����U  `�Some_stuffs_Some_stuffs_ �U  ����U   ���U  ����U   ���U  -5� /   ).� /       Meeting     �F��U  @G��U  �GSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �K��U  `V� /   {V� /       Some_stuffs `?��U  �?��U  `@Some_stuffs_Some_stuffs_ �U   C��U  �C��U  `D��U  �D��U  ��� /   ��� /       Some_stuffs �F��U  @G��U  �GSome_stuffs_Some_stuffs_ �U  PJ��U  �J��U  pK��U  �K��U  AЕ /   �ѕ /       Birthday    pc��U   d��U  �djustforfun_justforfun_ _ �U  �g��U   h��U  �h��U  0i��U  �� /   �� /      Some_stuffs �i��U  `j��U   kThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   p��U  �� /   a� /      Meeting     ���U  0��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `��U  -�� /   Ւ� /       Some_stuffs `?��U  �?��U  `@Some_stuffs_Some_stuffs_ �U   C��U  �C��U  `D��U  �D��U  ��� /   ɳ� /       Birthday    ����U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U   ݖ /   ݖ /       Birthday U  �u��U  `v��U   wThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   {��U  �� /   � /       Birthday    �� ��U  p� ��U  0� Some_stuffs_Some_stuffs_ �U  0� ��U   � ��U  �� ��U  �� ��U  �+� /   �+� /      Some_stuffs �
��U  ���U  �"justforfun_justforfun_ ��U   ��U  ���U   ��U  ���U  1R� /   rW� /      Workout     �� ��U  P� ��U  �� Some_stuffs_Some_stuffs_ �U  �� ��U  �� ��U   � ��U  �� ��U  � /   �~� /       Meeting     � ��U  �� ��U  �� justforfun_justforfun_  ��U  P� ��U  @� ��U  0� ��U  �� ��U  㡗 /   ʢ� /       Meeting     ����U   ���U  ��This_stuffs_This_stuffs_ �U   ���U  ����U  `���U   ���U  oŗ /   �˗ /       Appointment ����U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  � /   5� /      Workout      v��U  �v��U  `wSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  �{��U  N?� /   ><� /       Meeting     0[��U  �[��U  p\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  pa��U  �� /   <� /       Some_stuffs `���U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  X� /   �� /       Some_stuffs @� ��U   � ��U  �� Some_stuffs_Some_stuffs_ �U   ��U  ���U  @��U   ��U  �>� /   �9� /       Meeting ffs ���U  ����U  ��Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  �a� /   Re� /       Birthday     ���U  ����U  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �� /   `�� /       Some_stuffs Ѕ��U  ����U  @�justforfun_justforfun_ ��U  `���U  ����U  `���U  ����U  ű� /   볣 /       Meeting     �M��U  0N��U  �NSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �R��U  �ң /   �֣ /       Birthday    �� ��U  �� ��U   � This_stuffs_This_stuffs_ �U  `� ��U   � ��U  �� ��U  `� ��U  8�� /   ` � /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �(� /   �&� /      Appointment  � ��U  � ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p� ��U  >M� /   �M� /       Some_stuffs @���U  ���U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  9o� /   �q� /       Birthday    ����U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��� /   ��� /       Some_stuffs �� ��U  `� ��U   � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0� ��U  ��� /   �ä /       Some_stuffs                    justforfun_justforfun_ _Some_stuffs_Some_stuffs_             �� /   �� /      Appointment  5��U  �5��U   6This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   S��U  �� /   $� /       Some_stuffs ����U   ���U  p�This_stuffs_This_stuffs_ �U  p���U  ���U  ����U  @���U  8� /   58� /       Workout     �����U  `����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �\� /   �\� /      Birthday U  �3��U  �4��U   5Some_stuffs_Some_stuffs_ �U  @7��U   8��U  �8��U  @9��U  Z�� /   K�� /      Meeting     @����U  ����U  P��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��� /   ��� /       Workout     ����U  ����U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  Lҥ /   {ҥ /       Meeting     `>��U  �>��U  �?This_stuffs_This_stuffs_ �U  �B��U  `C��U   D��U  �D��U  ��� /   ��� /       Some_stuffs @���U   ���U  ��Some_stuffs_Some_stuffs_ �U   ���U  ����U  ����U  ���U  �!� /   �$� /       Workout     �� ��U  �� ��U  P� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   � ��U  �J� /   aC� /       Meeting      D��U  �D��U  �Ejustforfun_justforfun_ _ �U   H��U  �H��U  �U��U  pV��U  �m� /   �m� /      Meeting     @��U   ��U  �Some_stuffs_Some_stuffs_ �U  ���U  `	��U  �	��U  �
��U  ,�� /   A�� /       Meeting ent  g��U  �g��U  `hSome_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  �m��U  @� /   j� /      Meeting     @� ��U   � ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @ ��U  �� /   �� /      Meeting     ����U  p���U  �Some_stuffs_Some_stuffs_ �U   ���U  ����U  `���U   ���U  m3� /   �/� /       Birthday fs  >��U  �>��U   ?This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �B��U  �\� /   �\� /      Workout ffs ����U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  Џ��U  �*� /   X+� /       Some_stuffs `'��U  �'��U  �(Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p,��U  �V� /   �X� /      Birthday     J ��U  �J ��U  �N Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ` ��U  �|� /   �~� /       Some_stuffs �!��U  `"��U   #Some_stuffs_Some_stuffs_ �U  `%��U   &��U  �&��U   '��U  �� /   ��� /       Some_stuffs  G��U  �G��U   HSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   L��U  |ǲ /   �ǲ /      Some_stuffs � ��U  � ��U  � justforfun_justforfun_  ��U  0 ��U  � ��U  � ��U  � ��U  �� /   ;�� /       Birthday nt P� ��U  � ��U  �� Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  @� ��U  �� /   �� /       Meeting  fs �P��U  `Q��U   RThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �W��U  
h� /   �k� /       Some_stuffs ����U  ����U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  퍳 /   Y�� /       Some_stuffs                    This_stuffs_This_stuffs_                                     ŵ� /   ��� /      Meeting     PE��U  �E��U  �Fjustforfun_justforfun_ ��U   I��U  �I��U  PJ��U  �J��U  Uٳ /   �ܳ /       Workout ffs ����U  P���U  �This_stuffs_This_stuffs_ �U  ����U  ����U  P���U  ����U  �� /   � /       Some_stuffs  ���U  ����U  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  �-� /   �*� /       Meeting     ���U   ��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  N� /   VQ� /       Meeting      &��U  �&��U  `'justforfun_justforfun_ ��U  �)��U  P*��U  �*��U  p+��U  �z� /   �w� /      Some_stuffs  :��U  �:��U  �#This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p(��U  j�� /   ��� /       Some_stuffs P���U  У��U  ��justforfun_justforfun_ ��U  ����U  @���U  ����U  ����U  �Ǵ /   aǴ /       Birthday    p���U  0 ��U  � Some_stuffs_Some_stuffs_ �U  ���U  `��U  ���U  ���U  �� /   g� /      Some_stuffs ���U   ��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @��U  � /   u� /      Appointment  ���U  ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �7� /   �7� /      Meeting      ���U  ����U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  e� /   0e� /       Meeting     `� ��U   � ��U  �� justforfun_justforfun_  ��U  �� ��U  `� ��U  p� ��U  �� ��U  .�� /   ��� /       Appointment ���U   	��U  �	justforfun_justforfun_ _ �U  ���U  @��U   ��U  ���U  &�� /   ��� /       Some_stuffs �����U  @����U  ���Some_stuffs_Some_stuffs_ �U  �����U  P����U  �����U  @����U  ZԵ /   m۵ /       Birthday nt p,��U  �,��U  p-Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  p1��U  � /   F� /      Birthday nt 0b��U  �b��U  pcSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   h��U  �"� /   b(� /       Appointment ����U  p���U  ��This_stuffs_This_stuffs_ �U  @���U   ���U  ����U   ���U  DL� /   \L� /      Workout     ����U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `���U  �p� /   �s� /       Appointment ���U   ���U  ��justforfun_justforfun_ ��U  `���U   ���U  ����U  ����U  <�� /   ��� /       Meeting     pK��U  �K��U  pLThis_stuffs_This_stuffs_ �U  �N��U  pO��U  �O��U  pP��U  ��� /   �¶ /       Birthday     ���U  ����U  @�This_stuffs_This_stuffs_ �U  ����U  @���U   ���U  ����U  f7 &/   '7 &/       Birthday    @��U  ���U  @justforfun_justforfun_ ��U  `��U  ���U  ���U  	��U  ?_ &/   �_ &/       Some_stuffs ����U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  q� &/   � &/       Birthday nt ����U   ���U  �justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  `���U  � &/   �� &/       Some_stuffs �|��U  `}��U  ��Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  �� &/   � &/       Meeting      ���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  0� &/   I� &/      Workout �U  0O��U  �O��U  0PThis_stuffs_This_stuffs_ �U  `R��U  �R��U  `S��U  �S��U  $&/   6$&/      Meeting ent �� ��U  p� ��U  0� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  ,K&/   LK&/      Birthday    �U��U  pV��U  �IThis_stuffs_This_stuffs_ �U  �L��U  `M��U   N��U  �N��U  �n&/   il&/       Birthday     ��U  ���U  �	This_stuffs_This_stuffs_ �U  �"��U  @#��U  ���U  `��U  ��&/   ��&/       Workout ffs �$��U  �%��U  P&This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U   +��U  2�&/   x�&/       Appointment ����U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  L�&/   n�&/       Meeting                        This_stuffs_This_stuffs_                                     2
&/   �	&/       Some_stuffs �h��U  0i��U  �iSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `m��U  x0&/   �0&/      Workout                        This_stuffs_This_stuffs_                                     9\&/   �V&/       Appointment p/��U  00��U  �0This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  �5��U  5~&/   v�&/      Appointment ���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  8�&/   c�&/       Some_stuffs p+��U  �+��U  p,This_stuffs_This_stuffs_ �U  �.��U  p/��U  �/��U  p0��U  (�&/   3�&/      Birthday    �Y��U  �Z��U  0[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �_��U  X�&/   }�&/       Meeting     � ��U  �� ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  �&/   i&/       Some_stuffs 0,��U  �,��U  p-This_stuffs_This_stuffs_ �U  �/��U  �0��U  `1��U   2��U  �F&/   2G&/       Workout     P&��U  �1��U  �'This_stuffs_This_stuffs_ �U  `*��U   +��U  �+��U  �,��U  �h&/   �f&/       Meeting                        Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_             D�&/   |�&/       Appointment Pg��U  �g��U  p�justforfun_justforfun_ ��U   j��U  �j��U  `k��U  �k��U  4�&/   5�&/      Birthday fs ���U  ����U  `�This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U   ���U  �&/   �&/       Some_stuffs ����U  ����U  P�This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U   ��U  �2&/   �/&/      Appointment @� ��U   � ��U  �� This_stuffs_This_stuffs_ �U  � ��U  �� ��U  �� ��U  P� ��U  AW&/   fS&/       Workout     ���U  й��U  P�justforfun_justforfun_ ��U  ���U  н��U  P���U  ���U  ��&/   �&/      Workout     P����U  ����U  P��Some_stuffs_Some_stuffs_ �U  P����U  ����U  �����U  @����U  ��&/   ��&/       Some_stuffs �(��U  p)��U  �)justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  0.��U  �v&/   �|&/       Workout �U   &��U  �&��U  `'Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p+��U  %�&/   '�&/       Appointment `S��U   T��U  �TThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �Z��U  ��&/   ��&/       Some_stuffs p-��U  0.��U  �.justforfun_justforfun_ _ �U  `1��U   2��U  �2��U  @3��U  ��&/   ��&/      Meeting ffs ���U   ���U  ��This_stuffs_This_stuffs_ �U  `���U   ���U  ����U  ����U  �&/   �&/       Appointment ���U  ����U  0�justforfun_justforfun_ ��U  p���U  ����U  ����U  0���U  �<&/   �9&/       Birthday    �T��U  0U��U  �USome_stuffs_Some_stuffs_ �U  �W��U  pX��U   Y��U  �Y��U  �d&/   u_&/       Some_stuffs P���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U  ����U  P���U  ����U  y�&/   ��&/      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �&/   Q�&/       Meeting     �}��U  @~��U   justforfun_justforfun_ ��U  @���U   ���U  ����U   ���U  "�&/   %�&/       Appointment ����U  P���U  �Some_stuffs_Some_stuffs_ �U  л��U  ����U  ���U  н��U   &/   4&/       Some_stuffs ���U  p���U  0�justforfun_justforfun_ _ �U  ���U  p���U  ���U  p���U  =+&/   �(&/      Birthday    о��U  P���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  �M&/   VO&/      Birthday    P���U  ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Л��U  0x&/   ]x&/       Workout      o��U  �o��U   pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Pt��U  r�&/   ��&/       Birthday    ���U  p��U  Some_stuffs_Some_stuffs_ �U  ���U  ��U  ���U  ��U  ��&/   �&/       Workout ffs �N��U  pO��U  �OSome_stuffs_Some_stuffs_ �U  �Q��U  �R��U  pS��U  0T��U  ��&/   B�&/      Birthday    ���U   ��U  �justforfun_justforfun_ ��U   ��U  ���U   ��U  ���U  �&/   �&/       Workout     ����U  @���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  l6&/   �6&/      Workout  U  pF��U  �F��U  pGThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  PK��U  �\&/   `&/       Birthday    PE��U  �E��U  �FThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �J��U  ��&/   �&/       Meeting     `��U  ���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  X�&/   ~�&/      Some_stuffs `O��U  �O��U  `PSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  �U��U  ��&/   �&/       Workout     p� ��U  �� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   � ��U  !�&/   ��&/       Workout     �����U  P����U  ���justforfun_justforfun_ ���U  �����U  ����U  �����U  �  ��U  }%&/   � &/      Birthday    ����U  @���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  xG&/   �G&/       Appointment ����U  p���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  �n&/   �n&/       Birthday U  �h��U  �i��U  jThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Pn��U  +�&/   �&/       Birthday    �u��U  `v��U   wSome_stuffs_Some_stuffs_ �U  �y��U   z��U  �z��U   {��U  <�&/   g�&/      Meeting     P����U  ����U  P��Some_stuffs_Some_stuffs_ �U  P����U  ����U  �����U  @����U  D�&/   d�&/      Appointment 0���U  ���U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �&/   -
&/       Meeting �U  p=��U  �=��U  p>Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `u��U  �/&/   �/&/      Appointment  H��U  �H��U  �USome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `M��U  �T&/   Y&/      Workout  U   ���U  ����U  `�justforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U  ����U  U�&/   ?�&/       Appointment pL��U  �L��U  �MThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  pQ��U  9�&/   u�&/      Meeting     ���U  p���U  0�This_stuffs_This_stuffs_ �U  ����U  p���U  0���U  ����U  t�&/   ��&/      Birthday    �]��U  p^��U  0_Some_stuffs_Some_stuffs_ �U  0b��U  �b��U  �c��U  Pd��U  ��&/   N�&/       Some_stuffs �m��U  Pn��U  oSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   s��U   &/   � &/      Some_stuffs ����U  0���U  ��This_stuffs_This_stuffs_ �U  И��U  ����U  P���U  ���U  �C &/   a@ &/       Birthday    ���U  б��U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ж��U  �i &/   1j &/      Appointment �0��U  �1��U  02This_stuffs_This_stuffs_ �U  �4��U  �5��U  06��U  �6��U  �� &/   ?� &/      Workout     0b��U  �b��U  �cSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  h��U  �� &/   t� &/       Appointment ���U  б��U  ��Some_stuffs_Some_stuffs_ �U  ���U  ����U  ���U  ж��U  J� &/   /� &/       Birthday fs ���U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  �!&/   � !&/       Birthday    ���U  ���U  pThis_stuffs_This_stuffs_ �U  0��U  ���U  ���U   '��U  V+!&/   �*!&/       Birthday    @��U  ���U  @justforfun_justforfun_ ��U  @��U  ���U  `��U  ���U  ,S!&/   6S!&/       Birthday    ����U  0���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  w!&/   )w!&/      Birthday    �7 ��U  �8 ��U  @< justforfun_justforfun_  ��U  pE ��U  0F ��U   J ��U  �J ��U   �!&/   "�!&/      Appointment                    This_stuffs_This_stuffs_                                     ]�!&/   7�!&/       Workout     P&��U  �1��U  �'Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �,��U  �"&/   �"&/       Birthday    `��U   ��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ?"&/   �?"&/       Birthday    0� ��U   � ��U  �� justforfun_justforfun_  ��U  �� ��U  �� ��U   � ��U  �� ��U  �h"&/   @a"&/       Birthday    �k��U  l��U  �lThis_stuffs_This_stuffs_ �U  o��U  �o��U  �~��U   ��U  ��"&/   �"&/      Birthday    @��U   ��U  �Some_stuffs_Some_stuffs_ �U  ���U  ���U  ���U  0��U  x�"&/   {�"&/      Some_stuffs  ��U  ���U  �BThis_stuffs_This_stuffs_ �U  �!��U  `"��U   #��U  �#��U  �"&/   ��"&/      Meeting     ����U  @���U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  �(#&/   r,#&/       Birthday U   0��U  �0��U   =Some_stuffs_Some_stuffs_ �U  �3��U  �4��U   5��U  �5��U  �S#&/   �S#&/      Some_stuffs                    Some_stuffs_Some_stuffs_                                     ��-&/   z�-&/       Meeting      ��U  ���U  �This_stuffs_This_stuffs_ �U  ���U  ���U  `��U   ��U  l$.&/   ~$.&/       Meeting ffs ����U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ��U  �O.&/   �M.&/       Workout ffs  ]��U  �]��U  @^justforfun_justforfun_ _ �U  �`��U  Pa��U  �a��U  Pb��U  �q.&/   Nn.&/      Appointment pi ��U  0j ��U  �n justforfun_justforfun_  ��U  �z ��U  �{ ��U  0� ��U  �� ��U  ��.&/   k�.&/       Some_stuffs `��U  ���U  `This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `��U  2�.&/   y�.&/       Some_stuffs ���U   ��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @��U  !�.&/   �.&/       Birthday                       Some_stuffs_Some_stuffs_                                     �/&/   �/&/      Workout      � ��U  �� ��U  �� Some_stuffs_Some_stuffs_ �U  �� ��U  p� ��U  �� ��U  P� ��U  !3/&/   3:/&/      Birthday    `r��U   s��U  �sThis_stuffs_This_stuffs_ �U   v��U  �v��U  `w��U  �w��U  �_/&/   ?Z/&/       Birthday    R��U  �R��U  SSome_stuffs_Some_stuffs_ �U  PU��U  �U��U  PV��U  �V��U  ń/&/   ��/&/       Some_stuffs �����U  �����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  ��/&/   ��/&/       Some_stuffs �x��U  `y��U  �yjustforfun_justforfun_ ��U  �|��U  `}��U  ����U  p���U  ��/&/   ��/&/      Appointment �����U  �����U  ���Some_stuffs_Some_stuffs_ �U  �����U  @����U  �����U  @����U  ��/&/   ��/&/       Appointment @���U   ���U  ��This_stuffs_This_stuffs_ �U  p���U  ���U  ����U   ���U  �!0&/   �!0&/      Some_stuffs ����U  ����U  @�Some_stuffs_Some_stuffs_ �U   ���U  ����U  @���U  ����U  �F0&/   �F0&/      Appointment P#��U  $��U  �$This_stuffs_This_stuffs_ �U  �'��U   (��U  �(��U  �)��U  |q0&/   �q0&/       Workout     �s��U  `t��U  �tSome_stuffs_Some_stuffs_ �U  `w��U  �w��U  �x��U  `y��U  "�0&/   >�0&/       Some_stuffs                    justforfun_justforfun_                                       �0&/   �0&/      Workout     �����U  @����U   ��Some_stuffs_Some_stuffs_ �U  �����U  �  ��U  � ��U  � ��U  =�0&/   ��0&/      Appointment �4��U  p5��U  �5This_stuffs_This_stuffs_ �U  �8��U  9��U  �9��U  :��U  ,1&/   @1&/       Birthday    `���U  ����U  `�justforfun_justforfun_ ��U  `���U   ���U  ����U  ����U  �V1&/   �V1&/      Appointment � ��U  � ��U  � This_stuffs_This_stuffs_ �U   ! ��U  �! ��U  P% ��U  & ��U  ^�1&/   ��1&/       Workout     R��U  �R��U  SThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �V��U  !�1&/   �1&/       Birthday nt ���U  н��U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ^�1&/   ��1&/       Meeting     �2��U  p3��U  �3This_stuffs_This_stuffs_ �U  p6��U  07��U  �7��U  08��U  ��1&/   ?�1&/       Birthday     ��U  ���U  @Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  2&/   �2&/      Some_stuffs м ��U  �� ��U  P� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  �?2&/   �G2&/       Some_stuffs `1��U   2��U  �2justforfun_justforfun_ ��U   5��U  �5��U   6��U  �6��U  g2&/   �l2&/       Appointment  ��U  � ��U  @!Some_stuffs_Some_stuffs_ �U  @#��U  �#��U  @$��U  �$��U  YB=&/   �>=&/       Some_stuffs `h��U   i��U  �iSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �n��U  �c=&/   He=&/      Meeting     Pf��U  �f��U  PgSome_stuffs_Some_stuffs_ �U   i��U  �i��U   j��U  �j��U  �=&/   �=&/      Appointment p���U  ���U  ��This_stuffs_This_stuffs_ �U  `���U   ���U  ����U  ����U  =�=&/   ��=&/      Appointment `9��U  �9��U  �:Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  `@��U  n�=&/   ��=&/       Some_stuffs �a��U  Pb��U  �bSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �f��U  �>&/   X>&/       Workout     ����U  ����U  �Some_stuffs_Some_stuffs_ �U  ����U  ����U  ���U  ����U  �+>&/   �+>&/       Birthday nt `���U  ����U  ��This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  �T>&/   U>&/       Workout     �s��U  Pt��U  �tSome_stuffs_Some_stuffs_ �U  0w��U  �w��U  px��U  �x��U  �{>&/   �y>&/       Workout ffs `��U   ��U  �justforfun_justforfun_ ��U  `!��U  �!��U   :��U  �:��U  ��>&/   t�>&/       Workout     ����U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  ��>&/   ��>&/       Appointment P���U  П��U  ��justforfun_justforfun_ ��U  ����U  0���U  ����U  0���U  ��>&/   ��>&/       Workout     0� ��U  �� ��U  �� This_stuffs_This_stuffs_ �U  �� ��U  �� ��U  @� ��U   � ��U  �?&/   -?&/       Some_stuffs  ��U  ���U   This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  �7?&/   �7?&/       Meeting      N��U  �N��U  `OSome_stuffs_Some_stuffs_ �U   R��U  �R��U  `S��U   T��U  �a?&/   H^?&/       Meeting     P���U  ���U  ЮSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �?&/   �?&/      Workout     Ѕ��U  ����U  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  !�?&/   ��?&/      Some_stuffs �2��U  p3��U  �3This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  08��U  ��?&/   ��?&/       Some_stuffs ����U  `���U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  
@&/   }@&/       Some_stuffs `>��U  �>��U  �?Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �D��U  *@&/   0*@&/       Workout     ����U  ����U  `�This_stuffs_This_stuffs_ �U  `���U  ����U  ����U   ���U   J@&/   LJ@&/      Birthday    0����U  ����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p����U  �o@&/   r@&/       Meeting  U  ���U  0��U  �justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ���U  ��@&/   @&/       Appointment �� ��U  �� ��U  @� Some_stuffs_Some_stuffs_ �U   � ��U  �� ��U  �� ��U  @� ��U  ��@&/   9�@&/      Birthday    p���U  ����U  p�This_stuffs_This_stuffs_ �U  ���U  p���U  0���U  ���U  ��@&/   �@&/       Appointment P���U  ����U  p�justforfun_justforfun_ ��U  ����U  @���U  ����U  @���U  qA&/   �A&/       Meeting �U  �����U  �����U  ���justforfun_justforfun_ ���U  �����U  @����U  �����U  @����U  �5A&/   �5A&/       Appointment                    This_stuffs_This_stuffs_                                     �ZA&/   �\A&/       Workout �U  �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U  ہA&/   ��A&/       Appointment ����U  0���U  Иjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  P���U  "�A&/   ��A&/      Meeting     м ��U  �� ��U  P� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  ��A&/   ��A&/       Some_stuffs ����U  `���U   �justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  `���U  *�L&/   X�L&/       Workout     �[��U  @\��U   ]justforfun_justforfun_ ��U  �_��U  `��U  �`��U  Pa��U  p�L&/   ��L&/      Appointment �� ��U  @� ��U  �� Some_stuffs_Some_stuffs_ �U  � ��U  Щ ��U  �� ��U  � ��U  5�L&/   ��L&/       Workout  U  �����U  �����U  ���Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  @����U  Q�L&/   �L&/      Workout     ����U  p���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ?!M&/   �"M&/       Appointment �I��U  �J��U  `KThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �O��U  qBM&/   @IM&/       Some_stuffs p� ��U  �� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   � ��U  JjM&/   0pM&/       Some_stuffs ���U  `��U  This_stuffs_This_stuffs_ �U  @��U  ���U  @��U  ���U  M�M&/   ܖM&/       Workout     ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  P�M&/   �M&/       Meeting     �� ��U  p� ��U  0� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @� ��U  ��M&/   ��M&/       Some_stuffs �d��U  `e��U  �eThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `j��U  �N&/   �N&/       Appointment ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  1N&/   D1N&/      Birthday    �#��U  p$��U  0%This_stuffs_This_stuffs_ �U  �'��U  p(��U  �(��U  p)��U  M[N&/   IVN&/       Some_stuffs ����U  0���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p���U  �zN&/   {N&/      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��N&/   ȨN&/       Some_stuffs �����U  P����U  ���This_stuffs_This_stuffs_ �U  �����U  ����U  �����U  �  ��U  �N&/   @�N&/       Workout ent `_ ��U   ` ��U  `d Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �v ��U  pO&/   �O&/      Meeting     ���U  ���U  P Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �%��U  5@O&/   �CO&/      Appointment  %��U  �%��U   &This_stuffs_This_stuffs_ �U  �(��U  P)��U  �)��U  P*��U  �iO&/   _eO&/       Appointment �_��U  �`��U   aSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `e��U  J�O&/   �O&/      Appointment ����U   ���U  ��Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ����U  y�O&/   ݳO&/       Workout      ���U  ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ��O&/   ��O&/      Workout     p���U  0���U  ��This_stuffs_This_stuffs_ �U  ���U  Џ��U  P���U  ���U  LP&/   wP&/      Workout ffs ����U  p���U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �+P&/   �,P&/       Appointment �!��U  �"��U  P#Some_stuffs_Some_stuffs_ �U  P&��U  �1��U  �'��U   (��U  lRP&/   uRP&/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             FzP&/   �uP&/      Workout      ���U  ����U  @�This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  0���U  ��P&/   ��P&/       Workout     �� ��U  @ ��U   This_stuffs_This_stuffs_ �U  ���U  ���U  @��U   ��U  ��P&/   ��P&/       Workout ent �Z ��U  p[ ��U  `_ This_stuffs_This_stuffs_ �U  pi ��U  0j ��U  �n ��U  Po ��U  U�P&/   k�P&/       Workout ffs ����U  P���U  �justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ����U  ��[&/   x�[&/       Some_stuffs �����U  p����U  p��This_stuffs_This_stuffs_ �U  @����U  ����U  P����U  ����U  d�[&/   ��[&/      Meeting      � ��U  �� ��U  �� justforfun_justforfun_  ��U  �� ��U  `� ��U  �� ��U  �� ��U  �\&/   \&/      Meeting �U  м ��U  �� ��U  P� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U   5\&/   95\&/      Meeting �U   ��U  ���U   This_stuffs_This_stuffs_ �U  ���U   ��U  ���U  @��U  �a\&/   �a\&/       Some_stuffs  ���U  ����U   �This_stuffs_This_stuffs_ �U  @���U   ���U  ����U  @���U  B�\&/   ��\&/       Birthday    �����U  @����U  ���This_stuffs_This_stuffs_ �U  �����U  P����U  �����U  @����U  -�\&/    �\&/       Meeting     `� ��U   � ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  �\&/   �\&/       Workout ent PW��U   X��U  �XThis_stuffs_This_stuffs_ �U  �Z��U   [��U  �[��U  0\��U  � ]&/   D�\&/      Birthday     ]��U  �]��U  �^This_stuffs_This_stuffs_ �U   a��U  �a��U  `b��U   c��U  H#]&/   a#]&/      Birthday    @��U   ��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0��U  �L]&/   �H]&/       Appointment `���U  ����U  `�Some_stuffs_Some_stuffs_ �U  `���U   ���U  ����U  ����U  �p]&/   n]&/      Birthday    p���U  0���U  ��Some_stuffs_Some_stuffs_ �U  ����U  0���U  ����U  `���U  n�]&/   A�]&/       Some_stuffs ���U  ���U  pjustforfun_justforfun_ _ �U  0��U  ���U  ���U   '��U  ��]&/   ��]&/      Meeting     �����U  @����U  ���This_stuffs_This_stuffs_ �U  �����U  P����U  �����U  @����U  �]&/   )�]&/       Appointment `h��U   i��U  �iSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �n��U  �^&/   �^&/       Birthday                       justforfun_justforfun_ _                                     `2^&/   s2^&/      Some_stuffs Ю��U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  �W^&/   �W^&/       Birthday    0[��U  �[��U  p\This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  pa��U  �^&/   B�^&/       Birthday U  ����U  p���U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  M�^&/   ��^&/      Meeting �U  � ��U  � ��U  � Some_stuffs_Some_stuffs_ �U   ! ��U  �! ��U  P% ��U  & ��U  �^&/   ��^&/       Some_stuffs  |��U  �|��U  �}justforfun_justforfun_ ��U  @���U  ����U  @���U   ���U  ��^&/   �^&/       Workout     �@ ��U  �A ��U  pE This_stuffs_This_stuffs_ �U  �N ��U  �O ��U  �S ��U  �U ��U  �_&/   a"_&/       Birthday    P����U  ����U  P��Some_stuffs_Some_stuffs_ �U  P����U  ����U  �����U  @����U  �E_&/   �E_&/      Appointment �����U  `����U  ��justforfun_justforfun_ ���U  �����U  p����U  0����U  ����U  Ri_&/   !p_&/      Birthday    �*��U  p+��U  0,Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �0��U  �_&/   �_&/      Meeting     ���U  `��U   This_stuffs_This_stuffs_ �U  P��U  ���U  ���U  ���U  ȹ_&/   չ_&/      Workout     �P��U  `Q��U   Rjustforfun_justforfun_ ��U  �T��U  Pc��U  �V��U  �W��U  ��_&/   ��_&/       Workout      R��U  �R��U  `SSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0Y��U  �`&/   �`&/       Some_stuffs ����U  ���U  ��justforfun_justforfun_ ��U  д��U  P���U  е��U  ����U  Q1`&/   A0`&/       Workout     �� ��U  @� ��U   � This_stuffs_This_stuffs_ �U  �� ��U  p� ��U  �� ��U  P� ��U  �V`&/   =T`&/      Appointment @���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  0k&/   Zk&/      Meeting     `��U  ���U  `Some_stuffs_Some_stuffs_ �U  `��U  ���U  ���U  `��U  T1k&/   �1k&/       Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             _Qk&/   �Vk&/       Some_stuffs p/��U  00��U  �0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �5��U  �yk&/   �wk&/       Appointment P��U  ���U  �justforfun_justforfun_ ��U  ���U  ���U  p��U  ���U  e�k&/   D�k&/      Meeting     �O��U  P��U  �PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �T��U  ��k&/   ��k&/      Some_stuffs  ��U  ���U  @�Some_stuffs_Some_stuffs_ �U  ����U   ���U  ����U  @���U  ��k&/   4�k&/       Meeting     PE��U  �E��U  �FSome_stuffs_Some_stuffs_ �U   I��U  �I��U  PJ��U  �J��U  ^l&/   �l&/      Birthday nt `���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  �:l&/   �=l&/       Workout     `r��U   s��U  �sSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �w��U  (el&/   �jl&/       Meeting     ���U  ����U  �justforfun_justforfun_ ��U  ����U  ���U  ����U  ����U  T�l&/   Z�l&/      Some_stuffs �W��U  pX��U   YThis_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  �]��U  E�l&/   �l&/       Birthday    p8��U  �8��U  p9justforfun_justforfun_ _ �U  �;��U  p<��U  �<��U  p=��U  )�l&/   ��l&/       Appointment P���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  em&/   ��l&/       Workout     ����U  ����U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  t(m&/   �(m&/      Meeting     ���U   ��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `��U  �Mm&/   �Om&/      Meeting     �� ��U  @� ��U  �� Some_stuffs_Some_stuffs_ �U  � ��U  Щ ��U  �� ��U  � ��U  �sm&/   tm&/       Some_stuffs ����U  P���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  ��m&/   P�m&/       Meeting     ����U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  9�m&/   I�m&/       Workout      0��U  �0��U   =Some_stuffs_Some_stuffs_ �U  �3��U  �4��U   5��U  �5��U  �m&/   ��m&/      Birthday    @���U  ����U  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  Dn&/   Sn&/       Birthday    `'��U  �'��U  �(Some_stuffs_Some_stuffs_ �U  �*��U  p+��U  �+��U  p,��U  V8n&/   p<n&/       Workout     `r��U   s��U  �sSome_stuffs_Some_stuffs_ �U   v��U  �v��U  `w��U  �w��U  9^n&/   ~cn&/       Meeting     �� ��U  p� ��U  0� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  ��n&/   x�n&/       Some_stuffs п��U  P���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��n&/   �n&/       Meeting �U  ���U  `��U   justforfun_justforfun_ ��U  P��U  ���U  ���U  ���U  ��n&/   ��n&/       Meeting     px��U  �x��U  pyjustforfun_justforfun_ ��U  p{��U  �{��U  p|��U  0}��U  ��n&/   ��n&/       Workout     0� ��U  �� ��U  �� Some_stuffs_Some_stuffs_ �U  �� ��U  �� ��U  @� ��U   � ��U  'o&/   �#o&/       Meeting ffs �� ��U  �� ��U  P� Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U   � ��U  UKo&/   �Ho&/       Appointment �d��U  �e��U  PfThis_stuffs_This_stuffs_ �U  p���U  ����U   i��U  �i��U  �no&/   8so&/      Birthday    ����U   ���U  ��Some_stuffs_Some_stuffs_ �U  ����U  @���U  ����U  ����U  ]�o&/   B�o&/      Meeting     �	��U  �
��U  `justforfun_justforfun_ ��U   ��U  ���U  ���U  `��U  �Ez&/   �Ez&/       Some_stuffs `��U  ���U  �This_stuffs_This_stuffs_ �U  ���U   ��U  ���U  `��U  ��z&/   :�z&/       Some_stuffs �m��U  �n��U   oThis_stuffs_This_stuffs_ �U   q��U  �q��U   r��U  �r��U  νz&/   �z&/       Meeting     � ��U  � ��U  � justforfun_justforfun_  ��U  0 ��U  � ��U  � ��U  � ��U  ^
{&/   �{&/       Meeting ent �B��U  pC��U  ` This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  �$��U  m1{&/   7{&/       Birthday    �t��U  pu��U  0vjustforfun_justforfun_ ��U  px��U  �x��U  py��U  �y��U  �]{&/   y\{&/       Meeting       ��U  � ��U  `!Some_stuffs_Some_stuffs_ �U  �#��U  p$��U  0%��U  �%��U  6}{&/   �{&/      Meeting ffs ���U  ����U  P�justforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U   ���U  �{&/   |�{&/      Workout ffs ����U  ����U  @�justforfun_justforfun_ _ �U  ����U  @���U   ���U  ����U  t�{&/   u�{&/      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_              �{&/   G�{&/      Workout     �	��U   
��U  �
Some_stuffs_Some_stuffs_ �U  ���U  `��U   ��U  ���U   |&/   �|&/       Meeting     p=��U  �=��U  p>justforfun_justforfun_ ��U  �@��U  `A��U  �t��U  `u��U  %i|&/   j|&/       Birthday    �I��U  �J��U  `KThis_stuffs_This_stuffs_ �U  �M��U  �N��U  `O��U  �O��U  c�|&/   �|&/      Meeting     0��U  ���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  8�|&/   V�|&/      Appointment                    justforfun_justforfun_                                       a�|&/   ��|&/       Birthday    �'��U  p(��U  �(This_stuffs_This_stuffs_ �U  �*��U  p+��U  0,��U  �,��U  "}&/   }&/      Some_stuffs  ���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  H+}&/   _+}&/      Birthday    �����U  @����U  ���Some_stuffs_Some_stuffs_ �U  �����U  P����U  �����U  @����U  �Q}&/   #R}&/      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             Q}}&/   ��}&/      Meeting     �
��U  ���U  �"justforfun_justforfun_ ��U   ��U  ���U   ��U  ���U  )�}&/   H�}&/       Meeting     @���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  ��}&/   ��}&/       Workout     ����U  `���U  ��justforfun_justforfun_ ��U  `���U  ����U  ����U  `���U  �}&/   R�}&/       Birthday    ����U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U  �?~&/   �<~&/       Meeting      ���U  ����U  `�justforfun_justforfun_ _ �U  ����U  ����U  `���U   ���U  jc~&/   �c~&/       Some_stuffs �t��U  �u��U   vSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @z��U  |�~&/   ��~&/      Workout     ����U  @���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `���U  Ʒ~&/   l�~&/       Appointment  J ��U  �J ��U  �N Some_stuffs_Some_stuffs_ �U  �Z ��U  p[ ��U  `_ ��U   ` ��U  	��&/   ���&/       Appointment  ���U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  Ե�&/   �&/       Appointment  -��U  �-��U  �.This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   3��U  7؉&/   ۉ&/       Some_stuffs  ���U  ����U  @�This_stuffs_This_stuffs_ �U   ���U  ����U  `���U  ����U  P��&/   }��&/       Some_stuffs                    justforfun_justforfun_                                       v)�&/   �*�&/      Some_stuffs �@ ��U  �A ��U  pE This_stuffs_This_stuffs_ �U  �N ��U  �O ��U  �S ��U  �U ��U  �N�&/   �L�&/       Appointment � ��U  Щ ��U  �� This_stuffs_This_stuffs_ �U  P� ��U  p� ��U   � ��U  � ��U  �t�&/   �t�&/       Some_stuffs                    This_stuffs_This_stuffs_                                     ���&/   ˜�&/       Meeting      ���U  ����U  `�This_stuffs_This_stuffs_ �U  ����U  ����U  `���U  ����U  PŊ&/   ~Ŋ&/      Meeting     p\��U  0]��U  �]This_stuffs_This_stuffs_ �U  �`��U  pa��U  0b��U  �b��U  ��&/   (�&/       Some_stuffs ����U  ����U  `�justforfun_justforfun_ ��U  `���U  ����U  ����U   ���U  ��&/   n�&/      Meeting �U   � ��U  �� ��U  �� Some_stuffs_Some_stuffs_ �U  �� ��U  p� ��U  �� ��U  P� ��U  �:�&/   6:�&/       Meeting     `��U   ��U  �This_stuffs_This_stuffs_ �U  ���U  `��U  P��U  ���U  ���&/   ɂ�&/       Workout     ���U  @��U   This_stuffs_This_stuffs_ �U   ��U  ���U   ��U  0B��U  ��&/   ���&/       Meeting     P3 ��U  4 ��U  �7 justforfun_justforfun_  ��U  �@ ��U  �A ��U  pE ��U  0F ��U  $׋&/   G׋&/      Meeting ffs `D��U  �D��U  �ESome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  �J��U  ���&/   ���&/      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �&�&/   �%�&/       Workout     `!��U  �!��U   :This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �&��U  ,t�&/   It�&/       Appointment ���U  П��U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `���U  ғ�&/   V��&/       Appointment @n��U  �n��U  @ojustforfun_justforfun_ _ his_stuffs_This_stuffs_ �U  @t��U  ��&/   �&/      Birthday    �}��U  �~��U   Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  Ђ��U  2�&/   �8�&/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             V_�&/   �Z�&/      Some_stuffs  ��U  ���U   Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @��U  G��&/   脍&/       Appointment p� ��U  0� ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  Ǩ�&/   ���&/       Birthday    ����U  ����U  `�justforfun_justforfun_ _ �U   ���U  ����U  `���U   ���U  ��&/   ���&/       Meeting     `@��U   A��U  �AThis_stuffs_This_stuffs_ �U  `D��U  �D��U  �E��U  `F��U  X�&/   p�&/      Birthday    0����U  ����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p����U  �ј&/   �ɘ&/       Workout     ���U  @��U   This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ��U  ��&/   <��&/      Some_stuffs  -��U  �-��U  �.justforfun_justforfun_ ��U   =��U  �=��U  `2��U   3��U  (�&/   <�&/       Appointment ����U  `���U  �Some_stuffs_Some_stuffs_ �U  p���U  ����U  p���U  ����U  ]i�&/   �e�&/       Birthday     ���U  ����U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  �&/   ��&/      Birthday                       justforfun_justforfun_                                       2��&/   x��&/       Meeting ffs ����U  `���U   �justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  `���U  bݙ&/   ��&/       Meeting                        This_stuffs_This_stuffs_                                     ��&/   ��&/       Meeting     P���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  10�&/   M.�&/      Some_stuffs `O��U  �O��U  `PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �U��U  8P�&/   =P�&/      Appointment @� ��U   � ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  lz�&/   |�&/       Birthday    ����U  `���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  A��&/   p��&/      Some_stuffs �� ��U  @� ��U  �� justforfun_justforfun_  ��U  � ��U  Щ ��U  �� ��U  � ��U  �ƚ&/   �ƚ&/       Birthday    ����U  @���U  ��Some_stuffs_Some_stuffs_ �U  ����U  @���U   ���U  ����U  �&/   &�&/      Meeting     @���U  ����U  ��Some_stuffs_Some_stuffs_ �U   ���U  ����U  @���U  ����U  Y�&/   �&/       Meeting     ����U   ���U  ��justforfun_justforfun_ ��U  ����U  ���U  ����U  0���U  >�&/   G>�&/       Meeting      � ��U  �� ��U  @� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  �g�&/   �d�&/       Workout     `U��U  �U��U  �VThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   [��U  ���&/   ۍ�&/       Birthday    `d ��U   e ��U  pi This_stuffs_This_stuffs_ �U  �t ��U  �v ��U  �z ��U  �{ ��U  ���&/   ٳ�&/      Appointment �� ��U  P� ��U  �� This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  �� ��U  �ܛ&/   0֛&/       Some_stuffs �	��U  �
��U  `This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `��U  �&/   ���&/       Appointment `���U   ���U  ��This_stuffs_This_stuffs_ �U   ���U  ����U  `���U   ���U  _%�&/   �'�&/       Appointment `���U  ���U  ��justforfun_justforfun_ ��U  ���U  ����U  ���U  б��U  �O�&/   �O�&/      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ?��&/   ���&/       Birthday nt  w��U  �w��U  `xSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U   |��U  e&/   Fǜ&/       Birthday U  ���U  p��U  0This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  &�&/   ��&/       Birthday    p���U  ����U  p�Some_stuffs_Some_stuffs_ �U  ����U  `���U  ����U  `���U  n�&/   �&/       Meeting     `O��U  �O��U  �Pjustforfun_justforfun_ _ �U  `S��U   T��U  �T��U  Pc��U  �;�&/   =�&/       Workout     `U��U  �U��U  �VSome_stuffs_Some_stuffs_ �U  `Y��U  �Y��U  �Z��U   [��U  j�&/   |�&/       Some_stuffs ����U   ���U  ��justforfun_justforfun_ ��U  `���U   ���U  ����U  `���U  B5�&/   r6�&/       Appointment 0���U  ���U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  1Y�&/   _�&/      Some_stuffs �H��U  PI��U  Jjustforfun_justforfun_ _ �U  L��U  �L��U  PM��U  �M��U  l��&/   n��&/      Meeting     л��U  ����U  �This_stuffs_This_stuffs_ �U  ����U  ���U  ���U  ����U  ���&/   ���&/       Appointment  N��U  �N��U  `OThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   T��U  Ѩ&/   )Ѩ&/      Workout     � ��U  � ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  � ��U  o��&/   !��&/      Birthday    �����U  `����U  ��Some_stuffs_Some_stuffs_ �U  �����U  p����U  0����U  ����U  ��&/   ��&/       Workout     0� ��U  � ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  �H�&/   �H�&/      Birthday    07��U  �7��U  p8This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  p<��U  �n�&/   �n�&/      Appointment �� ��U  �� ��U   � justforfun_justforfun_  ��U  �� ��U  �� ��U  @� ��U   � ��U  K��&/   ��&/       Appointment �_��U  �`��U   aThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `e��U  |��&/   ���&/       Some_stuffs 0����U  ����U  ���justforfun_justforfun_ ���U   ����U  �����U  �����U  p����U  ��&/   {�&/       Meeting     `���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  �/�&/   �1�&/       Workout ent ���U  ���U  @This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  `	��U  Z�&/   �[�&/      Some_stuffs ���U  ���U  pSome_stuffs_Some_stuffs_ �U  p��U  ���U  ���U  p��U  ~�&/   L��&/       Appointment p��U  0��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  U��&/   �&/      Appointment �����U  @����U   ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  � ��U  �Ϫ&/   �˪&/       Meeting ffs P���U  Ђ��U  ��Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  ,�&/   [�&/       Appointment 0,��U  �,��U  p-Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   2��U  �?�&/   �G�&/       Meeting     �P��U  `Q��U   Rjustforfun_justforfun_ ��U  �T��U  Pc��U  �V��U  �W��U  Zj�&/   �i�&/       Meeting      ���U  ����U  `�This_stuffs_This_stuffs_ �U   ���U  ����U   ���U  ����U  I��&/   ���&/       Birthday    �!��U  �"��U  P#justforfun_justforfun_ _This_stuffs_This_stuffs_ �U   (��U  ���&/   ���&/       Appointment ���U   ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �$��U  9�&/   ��&/       Meeting �U  �����U  �����U  ���Some_stuffs_Some_stuffs_ �U  �����U  @����U  �����U  @����U  o�&/   �	�&/       Meeting      5��U  �5��U  �6This_stuffs_This_stuffs_ �U  `9��U  �9��U  �:��U  `;��U   0�&/   ;0�&/       Birthday    ���U  ���U  P This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �%��U  HV�&/   oV�&/      Appointment @� ��U   � ��U  �� Some_stuffs_Some_stuffs_ �U  � ��U  �� ��U  �� ��U  P� ��U  �z�&/   z�&/       Workout ffs �N��U  pO��U  �OSome_stuffs_Some_stuffs_ �U  �Q��U  �R��U  pS��U  0T��U  ؄�d�  ��/      Appointment �� ��U  p� ��U  0� This_stuffs_This_stuffs_ �U   � ��U  �� ��U  �� ��U  @� ��U  x#d�  ��/       Birthday U  `��U  ���U  �Some_stuffs_Some_stuffs_ �U  �	��U   
��U  �
��U  ���U  PLd�  84/      Appointment  -��U  �-��U  �.Some_stuffs_Some_stuffs_ �U   =��U  �=��U  `2��U   3��U  �)&d�  ��/       Meeting     `� ��U   � ��U  �� Some_stuffs_Some_stuffs_ �U  �� ��U  �� ��U  �� ��U  �� ��U  ��id�  �/      Some_stuffs   ��U  � ��U  `This_stuffs_This_stuffs_ �U  ���U  ���U  `��U  ���U  ���d�  H�/      Workout �U   A��U  �A��U  �BSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �G��U  �Zd�  ��/      Meeting �U  �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U  ȕd�  �/      Appointment p���U  0���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  8�Vd�  /�/      Some_stuffs �����U  �����U  ���Some_stuffs_Some_stuffs_ �U  �����U  @����U  �����U  @����U  ��N d�  pF/       Birthday                       justforfun_justforfun_                                       �(� d�  4m/      Workout     �� ��U  p� ��U  0� Some_stuffs_Some_stuffs_ �U   � ��U  �� ��U  �� ��U  @� ��U  x<�!d�  ]�/       Some_stuffs                    Some_stuffs_Some_stuffs_                                     �S�#d�  @/      Birthday     J ��U  �J ��U  �N justforfun_justforfun_  ��U  �Z ��U  p[ ��U  `_ ��U   ` ��U  (��Td�  $/      Meeting     ���U  `���U   �justforfun_justforfun_ ��U  ����U  `���U  ���U  ����U  x�Vd�  9�$/       Some_stuffs                    This_stuffs_This_stuffs_                                     �0�Vd�  :�$/      Some_stuffs ����U  @���U  ��justforfun_justforfun_ ��U  @���U  ����U  ����U  @���U  ��_Wd�  :%/      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��MYd�  @�%/      Appointment P��U  ���U  �This_stuffs_This_stuffs_ �U  ���U  ���U  p��U  ���U  ���]d�  �&/       Meeting     0���U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  8�^d�  ��&/      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �}bd�  h�'/       Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �\cd�  B�'/      Appointment �t��U  �u��U   vSome_stuffs_Some_stuffs_ �U  �x��U  `y��U  �y��U  �z��U  �J�d�  ��2/      Meeting     p� ��U  �� ��U   � justforfun_justforfun_  ��U   � ��U  �� ��U  @� ��U   � ��U  蛶�d�  G�3/      Appointment ����U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  П��U  �Ӛd�  ��4/       Workout     �� ��U  P� ��U  � justforfun_justforfun_  ��U  0� ��U  �� ��U  �� ��U  p� ��U  вz�d�  ��4/      Some_stuffs                    Some_stuffs_Some_stuffs_                                     �{@�d�  �5/      Birthday    0����U  ����U  ���This_stuffs_This_stuffs_ �U   ����U  �����U  �����U  p����U  ��՜d�  �A5/      Meeting �U  P� ��U  p� ��U   � justforfun_justforfun_ _ �U   � ��U  � ��U  �� ��U  �� ��U  X�x�d�  wg5/      Some_stuffs                    justforfun_justforfun_                                       ��/�d�  �5/      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��Ӟd�  Q�5/      Appointment �6��U   7��U  �7Some_stuffs_Some_stuffs_ �U  �:��U  `;��U   <��U  �<��U  ��/�d�  S	6/      Appointment p� ��U  �� ��U   � Some_stuffs_Some_stuffs_ �U   � ��U  �� ��U  @� ��U   � ��U  `٠d�  �06/      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             0�t�d�  �T6/       Birthday    p��U  0��U  �Some_stuffs_Some_stuffs_ �U  ���U  p��U  0��U  ���U  p^��d�  J�6/       Birthday    �m��U  Pn��U  oSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   s��U  `t �d�  �c7/      Some_stuffs �����U  `����U  ��This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  ����U  ��8�d�  /�B/       Appointment �� ��U  @� ��U  �� justforfun_justforfun_  ��U  � ��U  Щ ��U  �� ��U  � ��U  `���d�  .�C/      Birthday    ���U  ����U  P�Some_stuffs_Some_stuffs_ �U  ����U  ����U  ���U  ����U  ��6�d�  �C/       Workout     ���U  Џ��U  P�Some_stuffs_Some_stuffs_ �U  В��U  ����U  ���U  ����U  �n�d�  D7D/      Meeting     �����U  @����U   ��This_stuffs_This_stuffs_ �U  �����U  �  ��U  � ��U  � ��U  �I�d�  ܮD/      Some_stuffs �� ��U  P� ��U   � This_stuffs_This_stuffs_ �U  0� ��U  � ��U  �� ��U  p� ��U  ���d�  ��E/       Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��d�  ¨F/      Workout ent                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             p}�e�  DR/       Appointment                    Some_stuffs_Some_stuffs_                                     �(e�  lR/       Meeting �U  �=��U  �>��U  `?This_stuffs_This_stuffs_ �U  �A��U  �B��U   C��U  �C��U  ��Te�  )S/       Meeting     `� ��U   � ��U  �� justforfun_justforfun_  ��U  �� ��U  `� ��U  p� ��U  �� ��U  8�e�  [QS/      Birthday    �� ��U  p� ��U  0� justforfun_justforfun_  ��U  0� ��U   � ��U  �� ��U  �� ��U  : e�  ��S/       Some_stuffs @��U   ��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0��U  @� e�  ��S/       Some_stuffs pi ��U  0j ��U  �n Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  �A�$e�  E�T/      Some_stuffs `>��U  �>��U  �?This_stuffs_This_stuffs_ �U  �B��U  `C��U   D��U  �D��U  ~�%e�  C#U/       Birthday     J ��U  �J ��U  �N This_stuffs_This_stuffs_ �U  �Z ��U  p[ ��U  `_ ��U   ` ��U  ��&e�  �LU/       Some_stuffs � ��U  Ж ��U  �� This_stuffs_This_stuffs_ �U   � ��U  �� ��U  �� ��U  @� ��U  ��'e�  ��U/      Birthday    @� ��U   � ��U  �� justforfun_justforfun_ ��U   ��U  ���U  @��U   ��U  P�!)e�  0�U/       Some_stuffs �d��U  `e��U  �eSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `j��U  ��)e�  �V/      Appointment м ��U  �� ��U  P� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  `��Xe�  �a/      Birthday U  @��U   ��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0��U  X1iZe�  -`a/      Some_stuffs p� ��U  �� ��U   � Some_stuffs_Some_stuffs_ �U   � ��U  �� ��U  @� ��U   � ��U  �X\e�  Y�a/       Appointment �t ��U  �v ��U  �z justforfun_justforfun_  ��U  �� ��U  P� ��U   � ��U  �� ��U  h_e�  Krb/      Meeting ffs @7��U   8��U  �8This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   =��U  P�1be�  �/c/       Workout                        This_stuffs_This_stuffs_                                     ��/de�  ��c/      Meeting     P% ��U  & ��U  �) Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �8 ��U   �/fe�  �d/      Birthday    ���U  ���U  pThis_stuffs_This_stuffs_ �U  p��U  ���U  ���U  p��U  hZnge�  �gd/       Appointment �����U  @����U  ���This_stuffs_This_stuffs_ �U  �����U  P����U  �����U  @����U   ohe�  ,�d/       Workout     �� ��U  P� ��U   � justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  p� ��U  �!ie�  ��d/       Appointment 0<��U  �<��U  p=Some_stuffs_Some_stuffs_ �U  �?��U  0@��U  �@��U  `A��U  P�je�  �e/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             `lU�e�   p/       Some_stuffs �����U  �����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  ���e�  QPp/       Some_stuffs 0����U  ����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p����U  О��e�  \q/       Workout                        justforfun_justforfun_                                       ���e�  ��q/       Workout                        Some_stuffs_Some_stuffs_                                     Xѡe�  w�q/      Birthday nt ����U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  81�e�  �Kr/      Workout     �.��U  `/��U   0justforfun_justforfun_ ��U  `2��U   3��U  �3��U  �4��U  ��ƣe�  $sr/       Meeting      <��U  �<��U  `>justforfun_justforfun_ ��U   A��U  �A��U  �B��U  `C��U  ��ϥe�  Z�r/      Some_stuffs �� ��U  @� ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  � ��U  `�s�e�  �s/       Meeting     �t ��U  �v ��U  �z This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  8��e�  �6s/       Some_stuffs  ���U  ����U  `�This_stuffs_This_stuffs_ �U  ����U  ����U  `���U  ����U   ;��e�  ��s/      Appointment  Y��U  �Y��U  @ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �^��U  ȭ��e�  !D/      Some_stuffs @���U  ����U  ��This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U   ���U  ��R�e�  "=�/      Birthday    �t ��U  �v ��U  �z justforfun_justforfun_  ��U  �� ��U  P� ��U   � ��U  �� ��U  ����e�  8ځ/      Appointment `� ��U   � ��U  �� justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  �� ��U  hsC�e�  �'�/      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             8a��e�  �O�/       Workout ent �d��U  `e��U  �eThis_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  `j��U  Hi��e�  ʂ/      Birthday U  �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U  ��[f�  F��/      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             `�� f�  ���/       Birthday                       justforfun_justforfun_ _                                     �!f�  ���/       Meeting     �7 ��U  �8 ��U  @< Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �J ��U  ��#f�  ��/       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �$%f�  ʆ�/      Meeting     ���U  p��U  0This_stuffs_This_stuffs_ �U  P��U  ��U  ���U  ���U  ��'f�  ��/      Appointment �����U  @����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  �l�(f�  �p�/       Some_stuffs ���U  Л��U  ��This_stuffs_This_stuffs_ �U  ���U  П��U  ����U  @���U  �� *f�  ���/       Birthday    @����U   ����U  ���Some_stuffs_Some_stuffs_ �U  �����U  �����U  P����U   ����U  �e�+f�  �	�/      Some_stuffs p� ��U  0� ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  8#x-f�  �~�/       Appointment p� ��U  0� ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  X+cf�  ���/      Some_stuffs ���U  `��U   This_stuffs_This_stuffs_ �U  ���U  `��U  ���U  ���U  �8.ef�  �u�/      Some_stuffs  ��U  ���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0��U  pt�ff�  >ş/       Meeting ent  ��U  ���U   Some_stuffs_Some_stuffs_ �U  ���U   ��U  ���U   ��U  `c&gf�  *�/       Meeting                        This_stuffs_This_stuffs_                                     �r�hf�  f<�/       Meeting �U  `���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  �� if�  a�/      Workout     м ��U  �� ��U  P� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  �̴kf�  ���/       Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             @3hpf�  ��/       Some_stuffs  0��U  �0��U   =Some_stuffs_Some_stuffs_ �U  �3��U  �4��U   5��U  �5��U  �;��f�  	�/       Workout     `2��U   3��U  �3This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �8��U  �1#�f�  ^.�/      Birthday    ���U  й��U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  @���f�  ��/       Appointment �����U  p����U  p��This_stuffs_This_stuffs_ �U  @����U  ����U  P����U  ����U  0�Ѥf�  @E�/       Some_stuffs �+��U  p,��U  0-Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �1��U  X e�f�  �g�/       Some_stuffs �� ��U  P� ��U  �� Some_stuffs_Some_stuffs_ �U  �� ��U  �� ��U   � ��U  �� ��U  �½�f�  ѷ�/      Birthday nt �� ��U  �� ��U  0� justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  � ��U  `��f�  �-�/       Meeting     �����U  @����U   ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  � ��U  H�a�f�  /U�/       Some_stuffs ����U   ���U  �justforfun_justforfun_ ��U  `���U  ���U  ����U  `���U  ��f�  h��/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             H��f�  	��/      Workout     ���U  `��U   This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `��U  hж�f�  ��/       Birthday    ����U  ����U  p�This_stuffs_This_stuffs_ �U  P���U  ���U  Б��U  P���U  (�S�f�  7@�/       Workout     ����U  ����U  @�justforfun_justforfun_ ��U  ����U  ����U  @���U  ����U  h�f�  }۰/       Some_stuffs �^��U   _��U  �_Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `d��U  ؞<�f�  )�/       Birthday     A��U  �A��U  �BSome_stuffs_Some_stuffs_ �U  �E��U  `F��U   G��U  �G��U  �7��f�  v�/      Some_stuffs 0� ��U  �� ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   � ��U  �//�f�  �Q�/      Meeting ent ���U  p���U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �
�f�  d��/       Birthday     A��U  �A��U  �BThis_stuffs_This_stuffs_ �U  �E��U  `F��U   G��U  �G��U  8��f�  S;�/      Appointment                    This_stuffs_This_stuffs_                                     ح��f�  1Խ/       Workout     �� ��U  `� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0� ��U  (���f�  U#�/       Appointment �� ��U  @� ��U  `� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   � ��U  x���f�  �I�/      Birthday U  ���U  н��U  P�justforfun_justforfun_ ��U  ���U  ����U  ����U  ���U  ���f�  䚾/       Meeting ent p� ��U  �� ��U   � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   � ��U  x�H�f�  �/      Workout     0� ��U  �� ��U  �� This_stuffs_This_stuffs_ �U  �� ��U  @� ��U  � ��U  Ж ��U  P0�f�  xX�/       Birthday U  0����U  ����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p����U   �4�f�  �п/       Appointment  #��U  �#��U  `$Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  P(��U  ����f�  7l�/      Appointment �)��U  p*��U  �*Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p/��U  �
�f�  ���/      Meeting     ���U   ��U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  (Ƹ�f�  ���/      Workout      ��U  ���U  �BThis_stuffs_This_stuffs_ �U  �!��U  `"��U   #��U  �#��U  �d�}�  �T
 /      Birthday    0� ��U  � ��U  p� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0� ��U  x申}�  ) /      Appointment p� ��U  �� ��U   � Some_stuffs_Some_stuffs_ �U   � ��U  �� ��U  @� ��U   � ��U  ���}�  �S /       Appointment �� ��U  @� ��U  �� Some_stuffs_Some_stuffs_ �U  � ��U  Щ ��U  �� ��U  � ��U  {��}�  w /       Workout     @���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  X�P�}�  � /       Appointment �� ��U  �� ��U   � This_stuffs_This_stuffs_ �U  �� ��U  �� ��U  @� ��U   � ��U  h}�  �� /       Workout     ���U  ��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �#��U  P�G�}�   /      Workout     `_ ��U   ` ��U  `d This_stuffs_This_stuffs_ �U  �n ��U  Po ��U  �t ��U  �v ��U  �+�}�  �� /      Some_stuffs o��U  �o��U  �~This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `t��U  8
�}�  3p /       Appointment  � ��U  �� ��U  �� justforfun_justforfun_  ��U  �� ��U  p� ��U  �� ��U  P� ��U  p��}�  "� /      Appointment �^��U   _��U  �_justforfun_justforfun_ ��U  `b��U   c��U  �c��U  `d��U  ().�}�  W /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_              ���}�  �o /      Meeting     �� ��U  �� ��U  @� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @� ��U  !s�}�  � /       Birthday    � ��U  � ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  � ��U   ��}�  �� /      Some_stuffs  J ��U  �J ��U  �N Some_stuffs_Some_stuffs_ �U  �Z ��U  p[ ��U  `_ ��U   ` ��U  (u�}�  �� /       Workout ent  ���U  ����U  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �Q��}�  (? /      Some_stuffs p8��U  �8��U  p9This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p=��U  ��0~�  )) /       Appointment п ��U  �� ��U  P� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P� ��U  p�"2~�  �t) /       Workout �U  �� ��U  �� ��U  P� Some_stuffs_Some_stuffs_ �U  �� ��U  @� ��U  `� ��U   � ��U  �9�4~�  T* /       Birthday fs P���U  ���U  Юjustforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ���U  ��'6~�  yd* /       Appointment �� ��U  �� ��U  P� Some_stuffs_Some_stuffs_ �U  �� ��U  @� ��U  `� ��U   � ��U  �8~�  \�* /      Birthday    �(��U  p)��U  �)This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0.��U  h��8~�  �+ /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �Q<~�  E�+ /      Workout     P% ��U  & ��U  �) Some_stuffs_Some_stuffs_ �U  P3 ��U  4 ��U  �7 ��U  �8 ��U  ���<~�  v�+ /       Workout �U  0����U  ����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p����U  pT<=~�  V
, /       Meeting     p���U  0���U  ��This_stuffs_This_stuffs_ �U  ���U  Џ��U  P���U  ���U  `��=~�  7, /      Some_stuffs `?��U  �?��U  `@justforfun_justforfun_ _ �U   C��U  �C��U  `D��U  �D��U  ��?~�  ��, /       Meeting     �:��U  `;��U   <This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �A��U  �ŋ@~�  ��, /      Some_stuffs ����U  ���U  Юjustforfun_justforfun_ ��U  ����U  @���U  ���U  ����U  ��zB~�  �B- /       Some_stuffs �����U  @����U  ���Some_stuffs_Some_stuffs_ �U  �����U  P����U  �����U  @����U  �(�u~�  �,9 /      Some_stuffs ���U   ��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `��U  Mv~�  /R9 /       Appointment �� ��U  � ��U  Ы Some_stuffs_Some_stuffs_ �U   � ��U  � ��U  �� ��U  `� ��U  ��w~�  �}9 /       Birthday     ]��U  �]��U  @^This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Pb��U  p��y~�  �: /      Birthday                       justforfun_justforfun_                                       @JHz~�  b?: /      Appointment ���U  0��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `��U  `[�z~�  �c: /      Workout                        This_stuffs_This_stuffs_                                     pؚ}~�  R; /       Workout �U   ���U  ����U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U   ��~~�  hT; /       Workout     �� ��U  @� ��U  `� This_stuffs_This_stuffs_ �U   � ��U  �� ��U  �� ��U  `� ��U  �풁~�  ��; /       Meeting     �U��U  pV��U  �Ijustforfun_justforfun_ _ �U  �L��U  `M��U   N��U  �N��U  �[(�~�  �< /      Appointment  0��U  �0��U   =This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �5��U  ���~�  ��G /       Birthday    � ��U  @	 ��U  P Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  � ��U  �O�~�  8�G /       Meeting     ����U  @���U  ��justforfun_justforfun_ ��U  ����U   ���U  ����U  ����U  ���~�  �H /      Appointment � ��U  � ��U  � This_stuffs_This_stuffs_ �U   ! ��U  �! ��U  P% ��U  & ��U  @���~�  �JH /      Some_stuffs ����U  ����U  p�This_stuffs_This_stuffs_ �U  P���U  ���U  Б��U  P���U  ؋#�~�  iWI /       Meeting     �`��U  pa��U  0bThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �f��U  `!�~�  �-K /      Appointment ����U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  P�J�~�  ��V /       Some_stuffs  ���U  ����U  `�This_stuffs_This_stuffs_ �U  ����U  ����U  `���U   ���U  ���~�  ��V /       Workout     �� ��U  `� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  ����~�  �V /      Birthday    �Z ��U  p[ ��U  `_ Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  Po ��U  ����~�  �9W /       Some_stuffs ���U   ��U  �Some_stuffs_Some_stuffs_ �U   ��U  ���U   ��U  ���U  H1�~�  όW /       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ��#�~�  � X /       Appointment �����U  �����U  ���justforfun_justforfun_ ���U  �����U  @����U  �����U  @����U  �ܵ�~�  �X /       Some_stuffs                    Some_stuffs_Some_stuffs_                                     �U��~�  �Y /      Birthday U  ���U  0��U  �justforfun_justforfun_ ��U  `��U   ��U  ���U  `��U  Hzq�~�  �<Y /      Appointment �7 ��U  �8 ��U  @< Some_stuffs_Some_stuffs_ �U  pE ��U  0F ��U   J ��U  �J ��U  �SI�  ��Z /       Birthday U   � ��U  �� ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P� ��U  h��  k�Z /       Meeting     �:��U  0;��U  �;This_stuffs_This_stuffs_ �U  �=��U  p>��U  �>��U  p?��U  ����  ��Z /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             H.7�  �5f /       Some_stuffs ���U  ����U  оjustforfun_justforfun_ ��U  ���U  ����U  @���U  ����U  `Բ7�  rTf /      Some_stuffs �$��U  �%��U  P&This_stuffs_This_stuffs_ �U  �(��U  �)��U  `*��U   +��U  X�Z8�  �{f /       Appointment ���U   ��U  �Some_stuffs_Some_stuffs_ �U  `��U  ���U  ���U  `��U  @"9�  ��f /       Appointment                    Some_stuffs_Some_stuffs_                                     pEk:�  ��f /       Workout     0���U  ����U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �K;�  �g /       Birthday nt  v��U  �v��U  `wThis_stuffs_This_stuffs_ �U  �y��U  �z��U  `{��U  �{��U  x��;�  �?g /      Meeting �U  ����U  p���U  ��This_stuffs_This_stuffs_ �U  ����U  ����U  0���U  ����U  `{�>�  Xh /       Some_stuffs P� ��U  @� ��U  0� This_stuffs_This_stuffs_ �U  0� ��U  �� ��U  �� ��U  p� ��U  xڪ?�  ;/h /      Meeting      v��U  �v��U  `wSome_stuffs_Some_stuffs_ �U  �y��U  �z��U  `{��U  �{��U  ��GD�  Bi /      Appointment  A��U  �A��U  �BThis_stuffs_This_stuffs_ �U  �E��U  `F��U   G��U  �G��U  �9~G�  tj /       Workout     �:��U  `;��U   <This_stuffs_This_stuffs_ �U  �?��U  `@��U   A��U  �A��U  ���H�  EOj /      Appointment �����U  `����U  ��Some_stuffs_Some_stuffs_ �U  �����U  p����U  0����U  ����U  8��I�  �yj /      Appointment P����U  ����U  P��Some_stuffs_Some_stuffs_ �U  P����U  ����U  �����U  @����U  莝x�  pu /       Meeting     ����U   ���U  ��Some_stuffs_Some_stuffs_ �U  ����U  ���U  ����U  0���U  �hJy�  O�u /      Meeting     ���U  н��U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  ��	z�  ��u /       Some_stuffs �� ��U  `� ��U   � justforfun_justforfun_  ��U  0� ��U  � ��U  p� ��U  0� ��U  ���{�  �5v /       Appointment �����U  @����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  ���|�  1_v /       Appointment �� ��U  P� ��U  � Some_stuffs_Some_stuffs_ �U  0� ��U  �� ��U  �� ��U  p� ��U   ���  Fw /       Workout     �A��U  �B��U   CSome_stuffs_Some_stuffs_ �U  �E��U  `F��U  �F��U  �G��U  �얀�  ,Kw /      Appointment ���U  0��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `��U  ��|��  C�w /      Birthday                       justforfun_justforfun_                                       �ڃ�  �x /       Appointment �� ��U  p� ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  � ��U  H6��  �^x /       Birthday                       This_stuffs_This_stuffs_                                     ����  �|x /      Appointment 0����U  ����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p����U  �
q��  �y /      Some_stuffs � ��U  � ��U  � justforfun_justforfun_  ��U  0 ��U  � ��U  � ��U  � ��U  ���  e� /       Some_stuffs �� ��U  P� ��U  � This_stuffs_This_stuffs_ �U  � ��U  �� ��U  P� ��U  @� ��U  �z��  �ۄ /      Appointment 0%��U  �%��U  p&This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p*��U  Ȣ6��  ��� /      Some_stuffs ����U  P���U  �justforfun_justforfun_ ��U  л��U  ����U  ���U  н��U   
Ѿ�  �ƅ /      Birthday    ����U  ���U  ��This_stuffs_This_stuffs_ �U  ����U  ���U  ����U  P���U  �w���  ^�� /      Some_stuffs �����U  @����U   ��Some_stuffs_Some_stuffs_ �U  �����U  �  ��U  � ��U  � ��U  ����  �r� /       Meeting �U  �) ��U  P* ��U  �. Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   = ��U  �����  >�� /      Birthday    �t ��U  �v ��U  �z This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  PdU��   9� /      Some_stuffs ����U  ���U  �This_stuffs_This_stuffs_ �U  ����U  ����U  ���U  ����U  �����  �^� /      Meeting     г��U  ����U  �Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  й��U  �q���  �� /       Workout     P����U  ����U  P��Some_stuffs_Some_stuffs_ �U  P����U  ����U  �����U  @����U  X_j��  � /      Appointment �c��U  Pd��U  eThis_stuffs_This_stuffs_ �U  Pg��U  h��U  �h��U  �i��U  U���  �j� /      Meeting     ���U  ���U  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   '��U  � ��  75� /       Some_stuffs  ���U  ����U  ��Some_stuffs_Some_stuffs_ �U  @���U   ���U  ����U   ���U  �����  ã� /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             %���  UЕ /      Appointment �Z��U   [��U  �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0_��U  @DT��  �� /       Appointment  ���U  ����U   �Some_stuffs_Some_stuffs_ �U  ����U  `���U   ���U  ����U  �����  �� /       Meeting     �� ��U  P� ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p� ��U  X� ��  I�� /      Appointment �S ��U  �U ��U  �Z Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0j ��U  +���  � /      Appointment �t ��U  �v ��U  �z This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  ��5
��  XR� /       Appointment �t ��U  �v ��U  �z This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  P,�
��  � /      Birthday    �� ��U  @� ��U  `� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `� ��U  �h<��  �� /      Workout     �� ��U  �� ��U  @� This_stuffs_This_stuffs_ �U  �� ��U  @ ��U   ��U  ���U  Pq=��  �>� /       Meeting �U  p� ��U  �� ��U   � justforfun_justforfun_  ��U   � ��U  �� ��U  @� ��U   � ��U   �`?��  ��� /       Appointment о��U  P���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  HF�B��  Qo� /      Workout     �����U  @����U  ���Some_stuffs_Some_stuffs_ �U  �����U  P����U  �����U  @����U  ��I��  �!� /       Some_stuffs  � ��U  �� ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P� ��U  �Y�J��  �J� /      Meeting      0��U  �0��U   =Some_stuffs_Some_stuffs_ �U  �3��U  �4��U   5��U  �5��U  ���M��  �� /       Some_stuffs ����U  @���U  ��justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  ���U  ��qN��  �3� /      Workout     `���U  ���U  ��This_stuffs_This_stuffs_ �U  ���U  ����U  ���U  б��U  P��}��  �*� /       Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_              	N~��  W� /       Workout �U  � ��U  @	 ��U  P justforfun_justforfun_  ��U  � ��U  � ��U  � ��U  � ��U  p?���  P�� /      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             (�����  �� /      Appointment                    This_stuffs_This_stuffs_                                     訆���  #�� /       Workout     ���U  `��U   Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �g1���  ݵ� /       Appointment  � ��U  �� ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P� ��U  �m���  8� /       Meeting     @���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  0�����  �"� /       Birthday U  px��U  �x��U  pyThis_stuffs_This_stuffs_ �U  p{��U  �{��U  p|��U  0}��U  H�(J��  �� &/       Birthday nt ���U  ����U  @�justforfun_justforfun_ _This_stuffs_This_stuffs_ �U   ���U  �Y�J��  � &/      Birthday    �� ��U  P� ��U  � This_stuffs_This_stuffs_ �U  0� ��U  �� ��U  �� ��U  p� ��U   $R��  H\&/      Meeting                        This_stuffs_This_stuffs_                                     ��R��  g~&/       Birthday                       justforfun_justforfun_                                       (�V��  �h&/      Appointment  J ��U  �J ��U  �N Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ` ��U   �Z��  "3&/       Birthday    �t ��U  �v ��U  �z Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  0\�Z��  ^W&/      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ��q���  �v&/      Appointment `���U   ���U  �justforfun_justforfun_ ��U  ����U   ���U  ���U  `���U   � ���  V�&/       Meeting     �� ��U  @� ��U  `� justforfun_justforfun_  ��U  �� ��U  �� ��U  `� ��U   � ��U  �X���  �&/      Birthday    �t ��U  �v ��U  �z justforfun_justforfun_  ��U  �� ��U  P� ��U   � ��U  �� ��U   ����  ��&/       Some_stuffs �� ��U  `� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0� ��U  XVƑ��  a+&/       Some_stuffs                    justforfun_justforfun_                                       H"Z���  �M&/       Meeting ffs �����U  �����U  ���justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  @����U   8疗�  �\&/      Birthday    ���U  `���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  (�����  Y�&/      Workout     P����U  ����U  P��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  ��E���  �%&/       Appointment м ��U  �� ��U  P� justforfun_justforfun_  ��U  P� ��U  � ��U  �� ��U  �� ��U  p�dϗ�  ��&/      Meeting     �� ��U  `� ��U   � This_stuffs_This_stuffs_ �U  �� ��U  �� ��U   � ��U  �� ��U  �pЗ�  a�&/       Some_stuffs ����U  `���U  �justforfun_justforfun_ ��U  ���U  б��U  ����U  ���U  ���ї�  " &/       Meeting     ���U  н��U  P�Some_stuffs_Some_stuffs_ �U  ���U  ����U  ����U  ���U  x"�җ�  �C &/      Appointment ����U  `���U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �xGӗ�  j &/       Birthday    ���U   ��U  �Some_stuffs_Some_stuffs_ �U  `��U  ���U  ���U  `��U  ��ӗ�  Ќ &/       Meeting �U   0��U  �0��U   =This_stuffs_This_stuffs_ �U  �3��U  �4��U   5��U  �5��U  Ц)ٗ�  ��!&/      Birthday                       This_stuffs_This_stuffs_                                     �A�ۗ�  i"&/      Meeting     �� ��U  �� ��U  P� justforfun_justforfun_  ��U  �� ��U  @� ��U  `� ��U   � ��U  ��ܗ�  ��"&/       Meeting                        This_stuffs_This_stuffs_                                     pbߗ�  �(#&/      Meeting                        This_stuffs_This_stuffs_                                     �?���  �q.&/       Some_stuffs ����U  ���U  гjustforfun_justforfun_ ��U  ���U  ж��U  ����U  P���U  x���  K�.&/      Workout                        This_stuffs_This_stuffs_                                     P2���  B3/&/       Some_stuffs ���U  ���U    This_stuffs_This_stuffs_ �U   :��U  �:��U  �#��U  p$��U  P���  �_/&/       Some_stuffs �� ��U  p� ��U  0� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  � ��U  PE/��  ��/&/      Meeting �U  �� ��U  p� ��U  0� justforfun_justforfun_  ��U  @� ��U   � ��U  �� ��U  �� ��U  8�y��  ��/&/       Appointment � ��U  � ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  � ��U  x���  ��/&/       Birthday    P����U  ����U  P��This_stuffs_This_stuffs_ �U  P����U  ����U  �����U  @����U  �&��  E�0&/       Meeting �U  �����U  �����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @����U   IM��  $�1&/      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �RQ��  A2&/       Birthday                       justforfun_justforfun_                                       �9O��  �B=&/      Birthday U  �� ��U  p� ��U  0� This_stuffs_This_stuffs_ �U  0� ��U   � ��U  �� ��U  �� ��U  �Y�O��  �c=&/       Birthday     k��U  �k��U   mjustforfun_justforfun_ ��U  @o��U   p��U  �p��U  �q��U  ��Q��  e�=&/       Meeting     p���U  0���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  (�sR��  �>&/       Meeting     @� ��U   � ��U  �� justforfun_justforfun_ ��U   ��U  ���U  @��U   ��U  �J{T��  �{>&/       Workout     ���U  ����U  p�This_stuffs_This_stuffs_ �U  p���U  0���U  ����U  ����U  �ȺY��  U�?&/       Workout     ����U  ����U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  @�OZ��  ��?&/      Appointment � ��U  � ��U  � Some_stuffs_Some_stuffs_ �U   ! ��U  �! ��U  P% ��U  & ��U  `�2^��  ��@&/       Birthday    �� ��U  @� ��U  � justforfun_justforfun_  ��U  �� ��U  P� ��U   � ��U  �� ��U  ���^��  ��@&/      Some_stuffs Б��U  P���U  ВThis_stuffs_This_stuffs_ �U  P���U  ���U  ����U  P���U  �p�_��  �A&/       Workout      A��U  �A��U  �BSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �G��U  ��b��  ��A&/      Birthday    �7 ��U  �8 ��U  @< This_stuffs_This_stuffs_ �U  pE ��U  0F ��U   J ��U  �J ��U  ��
���  G�L&/       Birthday                       This_stuffs_This_stuffs_                                     ������  ��L&/       Meeting �U  п ��U  �� ��U  P� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P� ��U  ������  �BM&/       Workout �U  �P��U  `Q��U   RThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �W��U  PHU���  d�M&/      Appointment �� ��U  @� ��U  `� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   � ��U  �k����  ��M&/      Meeting �U   J ��U  �J ��U  �N Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ` ��U  0�I���  �N&/      Birthday                       Some_stuffs_Some_stuffs_                                     x˰���  m[N&/      Appointment �P��U  `Q��U   RSome_stuffs_Some_stuffs_ �U  �T��U  Pc��U  �V��U  �W��U  �����  c@O&/       Appointment �� ��U  @� ��U  �� Some_stuffs_Some_stuffs_ �U  � ��U  Щ ��U  �� ��U  � ��U   ~:���  �iO&/      Workout     ���U  `��U   Some_stuffs_Some_stuffs_ �U  P��U  ���U  ���U  ���U  0�����  ��O&/      Some_stuffs �l��U  Pm��U  �mThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �q��U  Ȇ5���  ��O&/       Appointment `{��U  �{��U  �|This_stuffs_This_stuffs_ �U  ���U   ���U  ����U  `���U  �|���  �+P&/       Some_stuffs `���U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  X6k���  �P&/      Appointment ����U  `���U   �justforfun_justforfun_ ��U  ����U  ����U  ���U  ����U   ����  ~�P&/      Meeting �U  �:��U  `;��U   <Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �A��U  `'R֘�  >�\&/      Workout �U  0����U  ����U  ���justforfun_justforfun_ ���U   ����U  �����U  �����U  p����U  8��ؘ�  �L]&/       Birthday    ���U  ����U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  hp�٘�  �p]&/       Birthday fs �\��U  0]��U  �]This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  �a��U  ��kۘ�  �]&/      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             p�5ܘ�  ^&/      Workout �U  �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U  ȅ�ޘ�  �^&/       Some_stuffs �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U  �&���  ��^&/       Some_stuffs �� ��U  @� ��U  �� Some_stuffs_Some_stuffs_ �U  � ��U  Щ ��U  �� ��U  � ��U  �����  �_&/      Workout                        Some_stuffs_Some_stuffs_                                     �����  �_&/      Some_stuffs                    justforfun_justforfun_                                       �=T��  g1`&/      Birthday                       justforfun_justforfun_                                       p<���  �V`&/       Workout                        justforfun_justforfun_                                       (����  �yk&/       Some_stuffs �����U  �����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @����U  `ł��  ��k&/       Some_stuffs `b��U   c��U  �cjustforfun_justforfun_ ��U  �e��U  `f��U   g��U  �g��U  @�/��  ��k&/       Birthday    ����U  ���U  Юjustforfun_justforfun_ ��U  ����U  @���U  ���U  ����U  �����  ��k&/      Appointment p� ��U  �� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   � ��U  P���  �:l&/       Meeting     �Q��U  �l��U  �Sjustforfun_justforfun_ ��U  �V��U  `W��U  �W��U  �X��U  (���  o�l&/       Workout                        This_stuffs_This_stuffs_                                     h+���  -�l&/      Some_stuffs `���U  ����U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U   b��  jm&/      Appointment �� ��U  � ��U  Ы This_stuffs_This_stuffs_ �U   � ��U  � ��U  �� ��U  `� ��U  �͸��  X�m&/      Some_stuffs                    Some_stuffs_Some_stuffs_                                     p�<"��  :^n&/      Meeting                        This_stuffs_This_stuffs_                                     �ʛ%��  'o&/       Birthday    ���U  П��U  ��This_stuffs_This_stuffs_ �U  `���U   ���U  ���U  `���U  ph8&��  �Ko&/       Workout ffs �d��U  �e��U  Pfjustforfun_justforfun_ _This_stuffs_This_stuffs_ �U  �i��U  ���&��  �no&/       Appointment ���U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  �'��  ��o&/       Meeting     @���U  ����U  ��Some_stuffs_Some_stuffs_ �U  `���U  ����U  `���U   ���U  �eU��  Fz&/      Appointment �7 ��U  �8 ��U  @< Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �J ��U  �#�V��  ��z&/      Some_stuffs  ��U  ���U  @Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  hwXY��  s1{&/      Birthday    `{��U  �{��U  �|This_stuffs_This_stuffs_ �U  ���U   ���U  ����U  `���U  �Z��  /^{&/      Workout                        This_stuffs_This_stuffs_                                      [�^��  Ji|&/      Birthday    �� ��U  p� ��U  0� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  `�`��  l�|&/      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �6c��  m}}&/       Meeting     �z ��U  �{ ��U  0� Some_stuffs_Some_stuffs_ �U   � ��U  �� ��U  �� ��U  @� ��U  P<�c��  N�}&/       Birthday    `� ��U   � ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `� ��U  ��=e��  6�}&/      Workout �U  �����U  �����U  ���justforfun_justforfun_ ���U  �����U  @����U  �����U  @����U  �{f��  @~&/      Some_stuffs  J ��U  �J ��U  �N Some_stuffs_Some_stuffs_ �U  �Z ��U  p[ ��U  `_ ��U   ` ��U  @����  ��&/       Meeting     �F��U  @G��U  �Gjustforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U  �K��U  8�I���  �N�&/      Some_stuffs                    Some_stuffs_Some_stuffs_                                     �郝��  ��&/       Appointment                    This_stuffs_This_stuffs_                                     x&9���  9��&/      Workout     � ��U  `� ��U  � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p� ��U  X�7���  '�&/       Some_stuffs �� ��U  P� ��U   � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `� ��U  �+����  2�&/      Birthday U  �� ��U  @� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P� ��U   <1ۙ�  ~i�&/      Appointment P% ��U  & ��U  �) Some_stuffs_Some_stuffs_ �U  P3 ��U  4 ��U  �7 ��U  �8 ��U  P5�ޙ�  :0�&/       Appointment �����U  @����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @����U  �aq���  N��&/       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ����  �ƚ&/      Birthday    � ��U  � ��U  � This_stuffs_This_stuffs_ �U   ! ��U  �! ��U  P% ��U  & ��U  ��y��  ^�&/       Some_stuffs ���U  p���U  0�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  X2��  1>�&/       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ����  �ܛ&/      Workout     �� ��U  @� ��U  `� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   � ��U  @(���  �&/      Birthday                       justforfun_justforfun_ _Some_stuffs_Some_stuffs_             ��_��  KY�&/       Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             h5���  ��&/       Appointment `K��U   L��U  �LThis_stuffs_This_stuffs_ �U  `O��U  �O��U  �P��U  `Q��U  ��D#��  �/�&/      Some_stuffs P#��U  $��U  �$Some_stuffs_Some_stuffs_ �U  �'��U   (��U  �(��U  �)��U  0��#��  <Z�&/       Appointment �� ��U  �� ��U  @� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  0�X%��  |��&/       Appointment  J ��U  �J ��U  �N justforfun_justforfun_ _ �U  �Z ��U  p[ ��U  `_ ��U   ` ��U  �c�'��  �?�&/       Meeting     �����U  @����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @����U  i')��  K��&/      Birthday U  �� ��U  p� ��U  0� Some_stuffs_Some_stuffs_ �U   � ��U  �� ��U  �� ��U  @� ��U  ��*��  K�&/      Some_stuffs                    justforfun_justforfun_                                       ��-��  �z�&/      Workout     0����U  ����U  ���This_stuffs_This_stuffs_ �U   ����U  �����U  �����U  p����U  �����O �/       Workout     `?��U  �?��U  `@This_stuffs_This_stuffs_ �U   C��U  �C��U  `D��U  �D��U  �3�p�O $p/      Workout      ���U  ����U  `�This_stuffs_This_stuffs_ �U   ���U  ����U    ��U  � ��U  �L�z�O 4/      Meeting     �����U  @����U   ��Some_stuffs_Some_stuffs_ �U  �����U  �  ��U  � ��U  � ��U  ����O �0/      Appointment �� ��U  p� ��U  0� This_stuffs_This_stuffs_ �U  0� ��U   � ��U  �� ��U  �� ��U  u��O è/       Birthday nt � ��U  �� ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  ��KI�O $/       Birthday                       justforfun_justforfun_                                       �V��O ��/       Workout �U  �7 ��U  �8 ��U  @< justforfun_justforfun_  ��U  pE ��U  0F ��U   J ��U  �J ��U  x۬�-�O W�#/      Birthday U  ����U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��,3.�O �#/       Meeting �U  ���U  p���U  0�justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  ����U  �i�1�O � &/       Workout     ���U  @��U   Some_stuffs_Some_stuffs_ �U  ���U  P��U   ��U  ���U  846�3�O �'/       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             _gEH�O �D3/      Birthday U  ���U  `��U   This_stuffs_This_stuffs_ �U  P��U  ���U  ���U  ���U  ���SI�O J�3/       Meeting                        justforfun_justforfun_ _                                      �đI�O �4/       Meeting     � ��U  � ��U  � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  � ��U  h�_�a�O �^B/       Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             Xi8�b�O C C/       Appointment �l��U  Pm��U  �mThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �q��U  0�{d�O ��C/      Appointment @r��U   s��U  �sjustforfun_justforfun_ ��U   v��U  �v��U   w��U  �w��U  H��d�O �D/       Meeting �U  �� ��U  `� ��U   � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0� ��U  8��~e�O ��D/      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ���Jf�O '�D/       Meeting     p� ��U  0� ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  �WJg�O �tE/       Workout                        This_stuffs_This_stuffs_                                      J�Rh�O 01F/       Some_stuffs 0���U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ���{�O �Q/      Birthday U  �����U  �����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  �X~�O ;S/      Meeting �U  ����U  `���U  �Some_stuffs_Some_stuffs_ �U  ���U  б��U  ����U  ���U  (on���O �!b/      Appointment �����U  `����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��'z��O ��c/       Appointment                    justforfun_justforfun_                                       p��D��O >Ed/      Workout �U  �����U  @����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @����U  0�+��O >�p/      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_              �ַ��O T�p/       Birthday    0� ��U  � ��U  p� Some_stuffs_Some_stuffs_ �U  0� ��U  � ��U  �� ��U  0� ��U  �#+y��O {aq/       Birthday U  �� ��U  �� ��U  @� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @� ��U  �z����O ��q/       Some_stuffs �. ��U  �/ ��U  P3 This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �A ��U  �i���O 
#r/      Some_stuffs  J ��U  �J ��U  �N justforfun_justforfun_  ��U  �Z ��U  p[ ��U  `_ ��U   ` ��U  Ȱ����O pt/       Appointment �P��U  `Q��U   RThis_stuffs_This_stuffs_ �U  �T��U  Pc��U  �V��U  �W��U  ݩ���O b�/       Workout                        justforfun_justforfun_                                       ��G��O �/       Some_stuffs @� ��U   � ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P� ��U  ��#��O ���/       Appointment �7 ��U  �8 ��U  @< This_stuffs_This_stuffs_ �U  pE ��U  0F ��U   J ��U  �J ��U  �դ7��O -�/      Appointment  J ��U  �J ��U  �N Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ` ��U  �DF���O �>�/       Workout     �� ��U  �� ��U   � This_stuffs_This_stuffs_ �U  �� ��U  �� ��U  @� ��U   � ��U  �(����O �c�/       Some_stuffs �����U  �����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  �Z� ��O ���/       Meeting      � ��U  �� ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Щ ��U  �7���O �!�/      Some_stuffs �����U  `����U  ��justforfun_justforfun_ ���U  �����U  p����U  0����U  ����U  XR)��O �N�/      Some_stuffs �P��U  `Q��U   RSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �W��U  �z����O �W�/      Appointment p� ��U  0� ��U  �� This_stuffs_This_stuffs_ �U  �� ��U  0� ��U  м ��U  �� ��U  ���z��O ��/      Birthday U  �� ��U  �� ��U  P� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   � ��U  x>h��O Β/      Appointment ���U  0��U  �justforfun_justforfun_ ��U  `��U   ��U  ���U  `��U  �1�+��O ��/       Appointment ���U  ����U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ����O ҈�/      Workout                        justforfun_justforfun_                                       �]���O �)�/       Birthday U  ���U  ����U  p�This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  X�O� �O ��/      Some_stuffs �����U  �����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @����U  0Ɣ�O ���/       Appointment ����U  p���U  �Some_stuffs_Some_stuffs_ �U   ���U  ����U  `���U   ���U  x�!�O w��/      Workout      J ��U  �J ��U  �N Some_stuffs_Some_stuffs_ �U  �Z ��U  p[ ��U  `_ ��U   ` ��U  �V�O �/       Some_stuffs `*��U   +��U  �+Some_stuffs_Some_stuffs_ �U  �.��U  `/��U   0��U  �0��U  @ٖ��O �߮/      Birthday                       Some_stuffs_Some_stuffs_                                     Hw�q�O щ�/       Appointment �� ��U  � ��U  Ы Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `� ��U  @E��2�O  ��/       Meeting     `� ��U   � ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  �ք4�O ���/       Some_stuffs  � ��U  �� ��U  �� This_stuffs_This_stuffs_ �U  �� ��U  p� ��U  �� ��U  P� ��U   ��M5�O D7�/      Some_stuffs @� ��U   � ��U  �� Some_stuffs_Some_stuffs_ �U  � ��U  �� ��U  �� ��U  P� ��U  ��P7�O �C�/       Meeting �U   � ��U  �� ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P� ��U  �R�-�O ��
 /       Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             h�1�2�O 5� /      Some_stuffs                    This_stuffs_This_stuffs_                                     H�p�F�O �� /       Some_stuffs ���U  Џ��U  P�This_stuffs_This_stuffs_ �U  В��U  ����U  ���U  ����U  ?$H�O �� /      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_              ���H�O � /       Some_stuffs  0��U  �0��U   =justforfun_justforfun_ ��U  �3��U  �4��U   5��U  �5��U  �od@J�O �� /       Workout     �?��U  `@��U   ASome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `F��U  (��J�O � /      Meeting     ����U  0���U  �This_stuffs_This_stuffs_ �U  ����U  @���U  ����U  ����U  �)�?K�O �| /       Workout      J ��U  �J ��U  �N This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ` ��U  ��6`�O Z�( /      Meeting �U  `���U  ����U  ��This_stuffs_This_stuffs_ �U  ����U   ���U  ����U  ����U  ��|a�O ��) /      Birthday U  �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U  ȇ�c�O q�* /       Meeting �U  �� ��U  �� ��U  P� justforfun_justforfun_  ��U  �� ��U  @� ��U  `� ��U   � ��U  8�}Lc�O ��* /       Meeting �U  `H��U   I��U  �IThis_stuffs_This_stuffs_ �U  �L��U  `M��U  �M��U  �N��U  @ݛd�O $+ /      Workout     м ��U  �� ��U  P� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  �Zf�O �X, /       Some_stuffs ���U  П��U  ��justforfun_justforfun_ ��U  `���U   ���U  ���U  `���U  ЩGog�O � - /       Birthday    `_ ��U   ` ��U  `d This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �v ��U  K{�O k�8 /       Birthday     � ��U  �� ��U  �� justforfun_justforfun_  ��U  �� ��U  p� ��U  �� ��U  P� ��U  �[{�O ��8 /       Appointment �|��U  `}��U  ��justforfun_justforfun_ ��U  ����U  `���U   ���U  ����U  8�6�O �*; /       Birthday    ����U  ���U  гjustforfun_justforfun_ ��U  ���U  ж��U  ����U  P���U  H����O Y�; /      Workout     ����U  p���U  �This_stuffs_This_stuffs_ �U   ���U  ����U  `���U   ���U  �=#:��O �; /       Some_stuffs �)��U  P*��U  �*justforfun_justforfun_ ��U  0-��U  �-��U  p.��U  �.��U  �0ܓ�O �[G /       Some_stuffs �z��U  �{��U   |This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��L��O ��H /       Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��3{��O ��H /      Birthday    ����U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  �G1���O ?�I /       Appointment @� ��U   � ��U  �� justforfun_justforfun_ ��U   ��U  ���U  @��U   ��U  P�S��O :�I /      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��V���O �J /       Appointment м ��U  �� ��U  P� Some_stuffs_Some_stuffs_ �U  P� ��U  � ��U  �� ��U  �� ��U  �ҵ̘�O $FJ /      Some_stuffs �7 ��U  �8 ��U  @< This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �J ��U  h���O �gJ /       Meeting ent P��U  ��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  $��U  x��V��O ��J /       Meeting     �� ��U  `� ��U   � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  �%$b��O ��K /      Meeting     �����U  `����U  ��Some_stuffs_Some_stuffs_ �U  �����U  p����U  0����U  ����U  ȥZ���O ɯW /       Workout �U  �����U  �����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U   b�ί�O ��W /       Some_stuffs ���U  ����U  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  x$w���O ��X /       Meeting     �����U  p����U  p��This_stuffs_This_stuffs_ �U  @����U  ����U  P����U  ����U  HӴݲ�O ��Y /       Appointment p� ��U  �� ��U   � Some_stuffs_Some_stuffs_ �U   � ��U  �� ��U  @� ��U   � ��U  @D�i��O ��Y /      Meeting     ���U  ���U  P This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �%��U  0:�7��O .vZ /      Birthday    �� ��U  P� ��U  � justforfun_justforfun_  ��U  0� ��U  �� ��U  �� ��U  p� ��U   m�$��O Hhg /       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ��7l��O x�g /       Workout �U  `Y��U  �Y��U  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   _��U  V���O kPh /       Workout                        justforfun_justforfun_                                       (�����O Mwh /       Meeting                        Some_stuffs_Some_stuffs_                                     0��>��O �h /       Appointment `K��U   L��U  �LSome_stuffs_Some_stuffs_ �U  `O��U  �O��U  �P��U  `Q��U  p����O v�h /       Birthday U  �.��U  p/��U  �/justforfun_justforfun_ ��U  �2��U  @3��U  �3��U  �4��U  h����O �i /       Birthday     � ��U  �� ��U  �� Some_stuffs_Some_stuffs_ �U  �� ��U  p� ��U  �� ��U  P� ��U  (����O gi /       Appointment `� ��U   � ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  pP��O n�i /      Birthday    `K��U   L��U  �LSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `Q��U  �:���O �Ku /       Appointment `���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U   {���O 0�w /      Appointment ���U  ���U  P This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �%��U  (����O M0x /      Workout �U  ����U  @���U  @Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �����O kgy /       Meeting �U  �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U   '���O �z� /       Some_stuffs                    Some_stuffs_Some_stuffs_                                     X����O �� /       Meeting     �� ��U  @� ��U  � justforfun_justforfun_  ��U  �� ��U  P� ��U   � ��U  �� ��U  (DJ���O ub� /       Meeting     0����U  ����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p����U  �~����O �)� /      Workout     �(��U  �)��U  `*Some_stuffs_Some_stuffs_ �U   -��U  �-��U  �.��U  `/��U   -�/ �O �P� /      Appointment �7 ��U  �8 ��U  @< Some_stuffs_Some_stuffs_ �U  pE ��U  0F ��U   J ��U  �J ��U  ��[�O �Г /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             H���O I�� /       Workout     �l��U  Pm��U  �mSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �q��U   Α��O ��� /       Meeting ent �2��U  @3��U  �3This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U   8��U  p��p�O n� /       Workout     �� ��U  @� ��U  `� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   � ��U   !u��O L?� /      Birthday nt pX��U  0Y��U  �YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p^��U  ���/�O �a� /      Some_stuffs �� ��U  � ��U  Ы Some_stuffs_Some_stuffs_ �U   � ��U  � ��U  �� ��U  `� ��U  ��(
1�O �(� /       Some_stuffs                    justforfun_justforfun_                                        QzH1�O lM� /      Meeting     ���U  ����U  �This_stuffs_This_stuffs_ �U  P���U  ����U  ����U  ���U  ��*S2�O �� /       Appointment �����U  `����U  ��Some_stuffs_Some_stuffs_ �U  �����U  p����U  0����U  ����U  ��N�2�O �� /       Birthday    �����U  `����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��2�O "8� /       Birthday    �� ��U  P� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p� ��U  ���X3�O f�� /       Appointment � ��U  � ��U  � This_stuffs_This_stuffs_ �U   ! ��U  �! ��U  P% ��U  & ��U  ��O4�O ��� /      Birthday                       Some_stuffs_Some_stuffs_                                     @Y=OI�O �|� /      Some_stuffs `d ��U   e ��U  pi justforfun_justforfun_  ��U  �t ��U  �v ��U  �z ��U  �{ ��U  h��J�O h� /       Birthday    0 ��U  � ��U  � Some_stuffs_Some_stuffs_ �U    ��U  � ��U   ! ��U  �! ��U  ��K�O �� /       Meeting     P����U  �����U  0��Some_stuffs_Some_stuffs_ �U  �����U  @����U  �����U  �����U  �8cL�O $N� /      Appointment                    justforfun_justforfun_                                        ��L�O �z� /       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_              -��L�O ��� /       Meeting �U  `{��U  �{��U  �|Some_stuffs_Some_stuffs_ �U  ���U   ���U  ����U  `���U  �:wN�O @�� /      Appointment  v��U  �v��U  `wThis_stuffs_This_stuffs_ �U  �y��U  �z��U  `{��U  �{��U  HJ��N�O 1�� /      Some_stuffs �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U  ��b�N�O �Ե /       Birthday    � ��U  � ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  � ��U   � P�O �p� /       Some_stuffs  � ��U  �� ��U  �� This_stuffs_This_stuffs_ �U  �� ��U  p� ��U  �� ��U  P� ��U  (���P�O ��� /       Some_stuffs                    Some_stuffs_Some_stuffs_                                     
�D�O �7 &/       Meeting     `� ��U   � ��U  �� Some_stuffs_Some_stuffs_ �U  �� ��U  `� ��U  p� ��U  �� ��U  h�p�F�O �n&/       Some_stuffs                    justforfun_justforfun_                                       �zDG�O ��&/       Birthday    �����U  @����U  ���Some_stuffs_Some_stuffs_ �U  �����U  P����U  �����U  @����U  8ϥ�G�O W�&/      Workout �U  �����U  �����U  ���Some_stuffs_Some_stuffs_ �U  �����U  @����U  �����U  @����U  x��H�O _
&/      Meeting �U  �����U  �����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @����U  8�1�I�O �&/      Meeting �U  �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U  �){T`�O �d&/      Appointment �� ��U  @� ��U  `� Some_stuffs_Some_stuffs_ �U  �� ��U  �� ��U  `� ��U   � ��U  �C��`�O '�&/      Appointment                    Some_stuffs_Some_stuffs_                                     ��a�O O�&/       Meeting     p\��U  0]��U  �]Some_stuffs_Some_stuffs_ �U  �`��U  pa��U  0b��U  �b��U  �[b�O ��&/      Appointment � ��U  � ��U  � Some_stuffs_Some_stuffs_ �U   ! ��U  �! ��U  P% ��U  & ��U   �U�b�O ��&/      Workout ent `���U   ���U  �Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  `���U   �.�b�O ��&/       Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �K@&c�O &/      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �;�c�O &/      Some_stuffs @< ��U   = ��U  �@ Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �O ��U  8!_%y�O �&/      Birthday nt @��U   ��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  8Q�y�O �T&/       Workout                        justforfun_justforfun_                                        춬z�O ��&/      Some_stuffs  J ��U  �J ��U  �N Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ` ��U   :|�O ̻ &/      Birthday     A��U  �A��U  �BSome_stuffs_Some_stuffs_ �U  �E��U  `F��U   G��U  �G��U  h�IB|�O M� &/      Birthday U  ���U  p��U  0This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  ���|�O [+!&/       Birthday    ����U  ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P���U   S&�~�O (?"&/      Some_stuffs �t ��U  �v ��U  �z This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  �� ��U  �L��O 9�"&/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             0w��O ��-&/       Workout      � ��U  �� ��U  �� Some_stuffs_Some_stuffs_ �U  �� ��U  p� ��U  �� ��U  P� ��U  `�� ��O �O.&/       Birthday U  0%��U  �%��U  p&justforfun_justforfun_ ��U  �(��U  p)��U  �)��U  p*��U  (��œ�O U�.&/       Workout      m��U  �m��U  @nThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   s��U  �e�Җ�O G�0&/       Appointment �����U  �����U  ���justforfun_justforfun_ ���U  �����U  @����U  �����U  @����U  �[i��O w�1&/      Meeting                        justforfun_justforfun_                                       �ʐ��O ��1&/       Workout �U  � ��U  � ��U  � Some_stuffs_Some_stuffs_ �U   ! ��U  �! ��U  P% ��U  & ��U  �S~X��O ��=&/       Meeting     �����U  @����U   ��This_stuffs_This_stuffs_ �U  �����U  �  ��U  � ��U  � ��U  ଺���O ��>&/      Meeting �U  �����U  �����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  �Ҟe��O �?&/       Appointment P����U  ����U  P��This_stuffs_This_stuffs_ �U  P����U  ����U  �����U  @����U  `�h���O 8?&/       Birthday    ���U  p��U  0Some_stuffs_Some_stuffs_ �U  P��U  ��U  ���U  ���U  8��O �a?&/      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��c.��O +�?&/       Workout     �	��U  �
��U  `Some_stuffs_Some_stuffs_ �U   ��U  ���U  ���U  `��U  hZ[���O -@&/      Meeting     p� ��U  �� ��U   � This_stuffs_This_stuffs_ �U   � ��U  �� ��U  @� ��U   � ��U  �����O �o@&/      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ��ĳ�O <�A&/       Birthday                       justforfun_justforfun_                                       xd,��O /�L&/      Meeting     `*��U   +��U  �+Some_stuffs_Some_stuffs_ �U  �.��U  `/��U   0��U  �0��U  (����O ejM&/       Meeting �U  `��U  ���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `��U  �olR��O `�O&/       Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �8����O _zP&/       Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �	i��O �P&/       Workout     P����U  ����U  P��justforfun_justforfun_ ���U  P����U  ����U  �����U  @����U  �CXF��O x�\&/      Some_stuffs `� ��U   � ��U  �� Some_stuffs_Some_stuffs_ �U  �� ��U  �� ��U  �� ��U  �� ��U  0����O � ]&/       Some_stuffs ���U  0��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `��U  �X���O ��]&/      Birthday    �s��U  @t��U  �tThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �x��U  �Y&���O W�^&/      Some_stuffs ���U  `��U   Some_stuffs_Some_stuffs_ �U  �
��U  ���U  �"��U  @#��U  �+�)��O Xi_&/       Birthday    ���U  ���U  P Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �%��U  P�f���O �l&/       Birthday    0����U  ����U  ���This_stuffs_This_stuffs_ �U   ����U  �����U  �����U  p����U  (����O -Nm&/       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �}�3��O ��m&/       Appointment �� ��U  p� ��U  0� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @� ��U  �����O B�m&/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��>��O k8n&/       Appointment �	��U  �
��U  `Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `��U  ���� �O  o&/       Birthday    �����U  `����U  ��This_stuffs_This_stuffs_ �U  �����U  p����U  0����U  ����U  8t�O ߽z&/      Appointment  5��U  �5��U  �6Some_stuffs_Some_stuffs_ �U  `9��U  �9��U  �:��U  `;��U  V���O j
{&/      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             h���O 5}{&/       Meeting                        This_stuffs_This_stuffs_                                     `�>U�O L}&/       Meeting     ����U  ����U  `�Some_stuffs_Some_stuffs_ �U  `���U  ����U  ����U   ���U  �H(0�O Է~&/       Some_stuffs `U��U  �U��U  �Vjustforfun_justforfun_ ��U  `Y��U  �Y��U  �Z��U   [��U  � e�.�O �)�&/       Birthday    В��U  ����U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  И��U  ���/�O �&/       Some_stuffs �Q��U  �l��U  �SSome_stuffs_Some_stuffs_ �U  �V��U  `W��U  �W��U  �X��U   ��a0�O ;�&/       Some_stuffs �����U  P����U  ���This_stuffs_This_stuffs_ �U  �����U  ����U  �����U  �  ��U  @Q�0�O ���&/       Some_stuffs 0� ��U  �� ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  �ۗ�2�O 㓌&/       Meeting �U  �� ��U  @� ��U  �� This_stuffs_This_stuffs_ �U  � ��U  Щ ��U  �� ��U  � ��U  xM24�O W_�&/       Appointment @����U   ����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ����U  ���H�O T��&/      Appointment �� ��U  P� ��U   � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `� ��U  ���*I�O zݙ&/      Meeting     `� ��U   � ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  P �rI�O �&/      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             (�1�K�O h�&/      Workout     @� ��U   � ��U  �� Some_stuffs_Some_stuffs_ �U   ��U  ���U  @��U   ��U  @�( L�O ���&/      Some_stuffs ����U  ���U  ЮSome_stuffs_Some_stuffs_ �U  ����U  @���U  ���U  ����U  x�F\N�O W�&/      Appointment `K��U   L��U  �LSome_stuffs_Some_stuffs_ �U  `O��U  �O��U  �P��U  `Q��U  @�ԜN�O p�&/      Meeting     `K��U   L��U  �LThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `Q��U  �!��N�O �;�&/      Appointment  J ��U  �J ��U  �N Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ` ��U  XΪ2a�O ��&/      Birthday    ���U  ���U  P justforfun_justforfun_ ��U  P#��U  $��U  �$��U  �%��U  ���ua�O G5�&/      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ����e�O �Ϫ&/      Appointment �V��U  `W��U  �WThis_stuffs_This_stuffs_ �U  �Z��U   [��U  �[��U  `\��U  ����f�O nj�&/      Some_stuffs �t ��U  �v ��U  �z Some_stuffs_Some_stuffs_ �U  �� ��U  P� ��U   � ��U  �� ��U  H�w2l��� /       Some_stuffs �t ��U  �v ��U  �z Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  ѫ�"MZ7�� /       Workout      A��U  �A��U  �BSome_stuffs_Some_stuffs_ �U  �E��U  `F��U   G��U  �G��U  ҫ�"MZ7�� /      Workout �U  `��U  ���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `��U  ӫ�"MZ7|� /       Appointment 0 ��U  � ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �! ��U  �-k9%dK�� /       Workout     ����U  `���U  ��justforfun_justforfun_ ��U  ����U  ����U  `���U  ����U  �-k9%dK� /       Appointment ����U  ����U  0�Some_stuffs_Some_stuffs_ �U  Ы��U  ����U  P���U  ���U  �-k9%dK^� /      Meeting     ����U  ���U  ��This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  P���U  ��
�/��%� /       Some_stuffs �����U  @����U   ��Some_stuffs_Some_stuffs_ �U  �����U  �  ��U  � ��U  � ��U  ��
�/��� /       Meeting     `b��U   c��U  �cjustforfun_justforfun_ ��U  �e��U  `f��U   g��U  �g��U  ��
�/��~� /       Workout ffs �~��U   ��U  �pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �u��U  !i�E���I /      Workout     �����U  @����U   ��Some_stuffs_Some_stuffs_ �U  �����U  �  ��U  � ��U  � ��U  "i�E���G /       Birthday U  ����U   ���U  p�Some_stuffs_Some_stuffs_ �U  p���U  ���U  ����U  @���U  #i�E��}D /       Workout ffs �� ��U  P� ��U  � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @� ��U  y��5j��� /       Some_stuffs �7 ��U  �8 ��U  @< This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �J ��U  z��5j��� /      Workout     p� ��U  0� ��U  �� This_stuffs_This_stuffs_ �U  �� ��U  0� ��U  м ��U  �� ��U  {��5j��� /       Meeting     �� ��U  @� ��U  `� This_stuffs_This_stuffs_ �U  �� ��U  �� ��U  `� ��U   � ��U  i��-V�)�H /      Some_stuffs @� ��U   � ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   � ��U  j��-V�)#�H /       Some_stuffs  ��U  ���U  0This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U   ��U  k��-V�)��H /       Meeting     ����U   ���U  ��Some_stuffs_Some_stuffs_ �U   ���U  ����U  `���U   ���U  )��{ϧ=�I /      Some_stuffs �t ��U  �v ��U  �z justforfun_justforfun_  ��U  �� ��U  P� ��U   � ��U  �� ��U  *��{ϧ=��I /       Appointment ���U  `��U   Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ���U  +��{ϧ=ڃI /       Meeting �U  @��U  ���U  `justforfun_justforfun_ ��U  �	��U  @
��U  �
��U  @��U  D�M���MZ /       Workout     `� ��U   � ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  D�M����KZ /       Workout     0����U  �����U  P��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �����U  D�M����NZ /       Appointment `��U   ��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �瞴03�[ /       Some_stuffs  � ��U  � ��U  �� justforfun_justforfun_  ��U  p� ��U  0� ��U  �� ��U  p� ��U  P��������&/       Workout     �����U  @����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  A!m�t�y /       Some_stuffs �� ��U  �� ��U  P� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   � ��U  B!m�tw�y /       Appointment �*��U  p+��U  0,This_stuffs_This_stuffs_ �U  �.��U  p/��U  �/��U  �0��U  C!m�tD�y /       Some_stuffs  ��U  ���U   This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  ���U  p��S�^N;� /       Meeting     P&��U  �1��U  �'This_stuffs_This_stuffs_ �U  `*��U   +��U  �+��U  �,��U  a�b;>��� /      Birthday    `���U   ���U  ��justforfun_justforfun_ ��U  `���U  ����U  ����U   ���U  b�b;>�x�� /       Meeting     �� ��U  �� ��U   � justforfun_justforfun_  ��U  `� ��U   � ��U  �� ��U  `� ��U  c�b;>�ı� /       Appointment `O��U  �O��U  `PSome_stuffs_Some_stuffs_ �U  �S��U  �T��U  `U��U  �U��U  �=x��S:�� /      Meeting      J ��U  �J ��U  �N justforfun_justforfun_  ��U  �Z ��U  p[ ��U  `_ ��U   ` ��U  �=x��S��� /       Appointment j��U  �j��U  �kSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �o��U  �=x��Sb�� /       Appointment �!��U  `"��U   #Some_stuffs_Some_stuffs_ �U  `%��U   &��U  �&��U   '��U  �ޯ�_�� /       Workout     В��U  ����U  �This_stuffs_This_stuffs_ �U  ����U  P���U  ���U  И��U  �ޯ�_e�� /       Meeting     `l��U  �l��U  �mSome_stuffs_Some_stuffs_ �U   p��U  �p��U   q��U  �q��U  �ޯ�_��� /       Meeting ffs 0v��U  �v��U  0wThis_stuffs_This_stuffs_ �U  py��U  �y��U  pz��U  �z��U  `��'�lٳ /      Some_stuffs `_ ��U   ` ��U  `d This_stuffs_This_stuffs_ �U  �n ��U  Po ��U  �t ��U  �v ��U  �Q��A�� /      Birthday    ����U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �Q��A�� /       Birthday fs ���U  `��U   Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @#��U  �Q��A?�� /       Appointment                    This_stuffs_This_stuffs_                                     9�d�|*�/       Appointment �]��U  p^��U  0_This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  Pd��U  !7�	&}*oo/       Meeting     `� ��U   � ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `� ��U  �����}*!/       Some_stuffs �� ��U  @� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P� ��U  Y�Un�}*_0/       Birthday    ����U   ���U  ��justforfun_justforfun_ ��U  ����U  @���U  ����U  ����U  �!��}*z�/      Workout     ����U  ���U  гSome_stuffs_Some_stuffs_ �U  ���U  ж��U  ����U  P���U  �"��%~*��/       Meeting     `� ��U   � ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  !T��B~*�/      Meeting     м ��U  �� ��U  P� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  �'���~*R�/       Appointment �� ��U  P� ��U  � Some_stuffs_Some_stuffs_ �U  0� ��U  �� ��U  �� ��U  p� ��U  �����*�#/       Meeting  U  P���U  ����U  P�justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ���U  �
�*��#/      Appointment 0� ��U  �� ��U  �� Some_stuffs_Some_stuffs_ �U  �� ��U  �� ��U  @� ��U   � ��U   ��ދ�*$�$/       Appointment `h��U   i��U  �iThis_stuffs_This_stuffs_ �U   m��U  �m��U  @n��U  �n��U  �6�x�*�=%/       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ��ar�*��%/       Some_stuffs p���U  ���U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0���U  9��Y(�*q'/      Appointment `� ��U   � ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  �L��s�*��'/       Some_stuffs 0����U  ����U  ���This_stuffs_This_stuffs_ �U   ����U  �����U  �����U  p����U  �h:"�*w!3/       Some_stuffs 0b��U  �b��U  �cSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  h��U  ���t9�*�F3/       Birthday U  �$��U  �%��U  P&This_stuffs_This_stuffs_ �U  �(��U  �)��U  `*��U   +��U  QE_$��*v�3/       Some_stuffs �Z��U   [��U  �[This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �`��U  �lL��*O
4/       Some_stuffs PN��U  O��U  �Ojustforfun_justforfun_ _This_stuffs_This_stuffs_ �U  �S��U  @H���*�T4/      Some_stuffs �t ��U  �v ��U  �z Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  �׋Y�*�z6/       Birthday                       This_stuffs_This_stuffs_                                     �җ|7�*�`B/      Some_stuffs ����U  ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  ,�w��*��B/       Meeting     ����U  P���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  1��>�*)�C/       Birthday    `?��U  �?��U  `@This_stuffs_This_stuffs_ �U   C��U  �C��U  `D��U  �D��U  	So�W�**D/      Workout     �� ��U  @� ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  � ��U  ��_(��*��D/       Some_stuffs �� ��U  `� ��U   � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0� ��U  9x��*@�D/      Meeting     �� ��U  @� ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  � ��U  xC(&�*/JE/       Meeting �U  `K��U   L��U  �Ljustforfun_justforfun_ ��U  `O��U  �O��U  �P��U  `Q��U  !wY(B�*�sE/       Some_stuffs   ��U  � ��U  `justforfun_justforfun_ ��U  ���U  ���U  `��U  ���U   ��u�*D�E/      Workout     0����U  ����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p����U  �$Hq��*��E/      Some_stuffs p� ��U  �� ��U   � Some_stuffs_Some_stuffs_ �U   � ��U  �� ��U  @� ��U   � ��U  ����*N6F/       Birthday    P���U  ����U  ��justforfun_justforfun_ ��U   ���U  ����U  ����U  @���U  �][Eל*�UF/       Meeting     `?��U  �?��U  `@Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �D��U  YHXj�*��Q/       Birthday U  �=��U  �>��U  `?Some_stuffs_Some_stuffs_ �U  �A��U  �B��U   C��U  �C��U  Hp+È�*i�Q/       Birthday nt  ���U  ����U  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  �#�N9�*.S/       Some_stuffs `2��U   3��U  �3justforfun_justforfun_ ��U  �6��U   7��U  �7��U  �8��U  P;n��*J~S/      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_             h�v���*�7a/       Meeting �U  �� ��U  � ��U  Ы Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `� ��U  itw�;�*#b/       Appointment 0��U  ���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  ࣴ���*\�b/       Some_stuffs ���U  `��U   justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ���U  hݴ��*M�b/       Workout      � ��U  �� ��U  �� This_stuffs_This_stuffs_ �U  @� ��U   � ��U  �� ��U  p� ��U  P��ӯ*Jc/      Workout �U  � ��U  � ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  & ��U  �Y�V�*��c/       Workout     �� ��U  �� ��U   � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   � ��U  �y�奰*nFd/       Meeting     ���U  ���U  `Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �!��U  @�ea��*�)p/       Birthday                       Some_stuffs_Some_stuffs_                                     ��и*ˠp/       Workout     �l��U  Pm��U  �mSome_stuffs_Some_stuffs_ �U  �~��U   ��U  �p��U  �q��U  ���*��p/       Appointment �~��U   ��U  �pSome_stuffs_Some_stuffs_ �U  �s��U  `t��U  �t��U  �u��U  �Ⱦ�R�*(`q/      Appointment ����U  ���U  дSome_stuffs_Some_stuffs_ �U  ���U  ����U  P���U   ���U  �X����*2�q/       Some_stuffs  A��U  �A��U  �BThis_stuffs_This_stuffs_ �U  �E��U  `F��U   G��U  �G��U  HCҗ��*��q/       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             Q4"�ҹ*�%r/       Appointment f��U  �f��U  PgSome_stuffs_Some_stuffs_ �U  j��U  �j��U  �k��U  l��U  (C�*"�*%�r/       Workout                        Some_stuffs_Some_stuffs_                                     he�@�*�Kt/       Meeting     ����U  @���U   �justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ���U  ��xX�*Yst/       Birthday    ���U  `	��U  �	Some_stuffs_Some_stuffs_ �U  ���U  `��U   ��U  ���U  P�3���*J�/       Some_stuffs @� ��U   � ��U  �� Some_stuffs_Some_stuffs_ �U   ��U  ���U  @��U   ��U  9�a��*T�/       Some_stuffs ����U  P���U  �Some_stuffs_Some_stuffs_ �U  ���U  Л��U  ����U  ���U  Y$���*\�/      Birthday                       This_stuffs_This_stuffs_                                     pI���*�1�/       Workout �U  �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U  �;�5j�*��/       Meeting �U  ����U  0���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  ��kԄ�*Xʀ/       Appointment �� ��U  p� ��U  0� This_stuffs_This_stuffs_ �U  0� ��U   � ��U  �� ��U  �� ��U  ���8!�*E��/      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             i��K��*��/       Appointment Ю��U  P���U  �Some_stuffs_Some_stuffs_ �U  ���U  ����U  `���U   ���U  !y �$�*�>�/       Some_stuffs  j��U  �j��U  `kSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �o��U  )A	=�*�e�/      Meeting      � ��U  �� ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  �)���*į�/       Appointment �@��U  �A��U  0BSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @G��U  P�	��*�֎/       Appointment ���U  ����U  P�This_stuffs_This_stuffs_ �U  P���U  ����U  ����U   ���U  IÅ�*�#�/       Workout     �����U  `����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  W���*�H�/       Appointment  5��U  �5��U   6This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   S��U  @��8�*(t�/       Birthday     � ��U  � ��U  �� Some_stuffs_Some_stuffs_ �U  p� ��U  0� ��U  �� ��U  p� ��U  	C!��*�X�/       Birthday    `� ��U   � ��U  �� This_stuffs_This_stuffs_ �U  �� ��U  `� ��U  p� ��U  �� ��U  �~֭�*Ъ�/       Workout ent `>��U  �>��U  �?justforfun_justforfun_ ��U  �B��U  `C��U   D��U  �D��U   7E���*d��/       Appointment                    justforfun_justforfun_                                       �/�p�*ɒ/       Meeting     �M��U  0N��U  �NSome_stuffs_Some_stuffs_ �U  �P��U  pQ��U  �Q��U  �R��U  ћ����*��/      Some_stuffs �� ��U  `� ��U  p� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U   1B�*�d�/       Some_stuffs �� ��U  @� ��U  `� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   � ��U  �Ҡ3�*���/       Birthday    0���U  Щ��U  ��Some_stuffs_Some_stuffs_ �U  P���U  ���U  Ю��U  ����U  1I����*w(�/       Appointment ����U  p���U  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �KR@5�*��/       Workout �U  ����U  @���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  8n�m��*筠/       Workout     �� ��U  �� ��U  @� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @� ��U  p�I �*.r�/      Birthday     ��U  ���U   Some_stuffs_Some_stuffs_ �U  ���U  `��U   ��U  ���U  qZ�S6�*ߣ�/      Appointment ���U  `��U   This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  �#�xh�*���/       Appointment �i��U  `j��U   kjustforfun_justforfun_ ��U  @n��U  �n��U  @o��U   p��U  �w���*
�/       Some_stuffs P ��U  !��U  �!This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �1��U  ����*�/       Some_stuffs �V��U  pW��U  �Wjustforfun_justforfun_ ��U  @Z��U   [��U  �[��U  @\��U  ��<��*��/       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ��ˎ8�*ճ�/       Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             X� m�*K�/       Appointment `� ��U   � ��U  �� This_stuffs_This_stuffs_ �U  �� ��U  `� ��U  p� ��U  �� ��U  ��]���*�p�/       Some_stuffs ���U  н��U  P�Some_stuffs_Some_stuffs_ �U  ���U  ����U  ����U  ���U  �}aN�*�/       Workout     0����U  ����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p����U  �3���*&��/       Some_stuffs  q��U  �q��U   rThis_stuffs_This_stuffs_ �U  `t��U  ���U  �u��U  `v��U  z�\��*���/       Meeting ffs �?��U  `@��U   ASome_stuffs_Some_stuffs_ �U   D��U  �D��U  �E��U  `F��U  !b����*A/�/       Some_stuffs �h��U  �i��U  jSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  Pn��U  O|n��*�H�/       Appointment  � ��U  �� ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P� ��U  �jt�m.Q~
 /       Workout     �� ��U  P� ��U   � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p� ��U  �l[�m.��
 /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��(~�m.k�
 /      Some_stuffs �� ��U  `� ��U   � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0� ��U  ��U^�m.[ /      Birthday    � ��U  � ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  � ��U   I��Gn.$� /       Some_stuffs �t ��U  �v ��U  �z This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  p_+ao.�9 /       Birthday    p� ��U  �� ��U   � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   � ��U  �o.� /       Meeting �U  � ��U  � ��U  � Some_stuffs_Some_stuffs_ �U  0 ��U  � ��U  � ��U  � ��U  ��B�o.R  /       Workout     @���U   ���U  ��This_stuffs_This_stuffs_ �U  p���U  ���U  ����U   ���U  p���p.R /       Workout      � ��U  �� ��U  �� Some_stuffs_Some_stuffs_ �U  �� ��U  p� ��U  �� ��U  P� ��U  	:;�w.@� /      Appointment ���U  `��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  � ��U  �O�)x.�~ /      Appointment 0����U  ����U  ���Some_stuffs_Some_stuffs_ �U   ����U  �����U  �����U  p����U  ���Cx.ȥ /       Birthday U  �� ��U  @� ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  � ��U  ���^x.2� /      Meeting     `���U  ����U  ��Some_stuffs_Some_stuffs_ �U   ���U  ����U  `���U  ����U  A4ľ�x.9! /       Meeting                        This_stuffs_This_stuffs_                                     9�5�y.t� /      Some_stuffs `!��U  �!��U   :Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �&��U  ��{�/y.� /       Workout     ���U  Л��U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U   %k�Dy.�+ /       Meeting     @����U   ����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ����U  iI�Wzy.�� /       Meeting     ���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  8�6��y.'� /      Meeting �U   A��U  �A��U  �BThis_stuffs_This_stuffs_ �U  �E��U  `F��U   G��U  �G��U  (�D�y.A /       Appointment 0����U  ����U  ���justforfun_justforfun_ ���U   ����U  �����U  �����U  p����U  �2��.z.8� /      Meeting      0��U  �0��U   =This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �5��U  �K����.�( /       Meeting     `� ��U   � ��U  �� justforfun_justforfun_  ��U  �� ��U  �� ��U  �� ��U  �� ��U  ���h*�.,�) /       Workout     ����U  @���U   �Some_stuffs_Some_stuffs_ �U  ����U  ����U  @���U   ���U  ���F�.��) /      Birthday    @o��U   p��U  �pSome_stuffs_Some_stuffs_ �U  �s��U  @t��U  �t��U  �u��U  ��u9Ƃ.��* /       Workout     �����U  `����U  ��Some_stuffs_Some_stuffs_ �U  �����U  p����U  0����U  ����U  y=ч߂.��* /       Some_stuffs �t��U  �u��U   vSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @z��U  �Kg�,�.$+ /       Workout      � ��U  �� ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P� ��U  �j����.�Z, /      Meeting ent �� ��U  �� ��U  @� justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  @� ��U  ��F(}�.�!- /       Workout       ��U  � ��U  `This_stuffs_This_stuffs_ �U  ���U  ���U  `��U  ���U  �i_Ë.:8 /      Workout     ���U  ����U  ��This_stuffs_This_stuffs_ �U  ���U  ����U  P���U  ����U  0��U�.��8 /       Appointment �� ��U  �� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   � ��U  Y��f)�.¶8 /      Workout �U  ���U  p���U  �justforfun_justforfun_ ��U  0���U  ���U  ����U  p���U  9�jkE�.��8 /      Birthday U   ��U  ���U  @�Some_stuffs_Some_stuffs_ �U  ����U   ���U  ����U  @���U  y$�Ǎ.".; /      Workout     �����U  @����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @����U  `�7���.�u; /      Some_stuffs                    justforfun_justforfun_                                       ɟ�N�.i�; /       Workout ffs ���U   ��U  ��justforfun_justforfun_ _ �U  ����U  @���U  ����U  p���U  �#:�,�.�; /      Appointment  5��U  �5��U   6Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   S��U  Q}�ؕ.X^G /       Birthday    ����U  ����U  @�justforfun_justforfun_ ��U  ����U  ����U  @���U  ����U  ������.��G /       Birthday     0��U  �0��U   =justforfun_justforfun_ ��U  �3��U  �4��U   5��U  �5��U  ������.K�H /      Meeting     �� ��U  p� ��U  0� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  �#
=ޖ.h�H /       Appointment ����U  `���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �=(��.Y
I /      Birthday                       Some_stuffs_Some_stuffs_                                     ���[�.שI /       Appointment  0��U  �0��U   =justforfun_justforfun_ ��U  �3��U  �4��U   5��U  �5��U  �1mw�.��I /       Some_stuffs �*��U  p+��U  0,Some_stuffs_Some_stuffs_ �U  �.��U  p/��U  �/��U  �0��U  ��_+��.�J /       Workout      � ��U  �� ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   � ��U  !C(Ɨ.-FJ /       Workout      J ��U  �J ��U  �N This_stuffs_This_stuffs_ �U  �Z ��U  p[ ��U  `_ ��U   ` ��U  ���{ܗ.�pJ /       Birthday    ���U  ���U  `This_stuffs_This_stuffs_ �U   ��U  ���U  �	��U   
��U  9c7
��.׏J /       Some_stuffs ����U   ���U  ��justforfun_justforfun_ ��U   ���U  ����U   ���U  ����U  �ogx�.�SK /       Workout �U  �� ��U  p� ��U  0� Some_stuffs_Some_stuffs_ �U  0� ��U   � ��U  �� ��U  �� ��U  �3v��.��K /       Some_stuffs �� ��U  p� ��U  0� This_stuffs_This_stuffs_ �U  0� ��U   � ��U  �� ��U  �� ��U  1!6~Ș.?�K /       Appointment  � ��U  �� ��U  �� Some_stuffs_Some_stuffs_ �U  �� ��U  p� ��U  �� ��U  P� ��U  Ik�	��.a�W /       Meeting     P� ��U  @� ��U  0� This_stuffs_This_stuffs_ �U  0� ��U  �� ��U  �� ��U  p� ��U  �-2à.��W /       Appointment `U��U  �U��U  �VSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   [��U   �!S�.`MX /       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             �?�\�.��X /       Meeting �U  ���U  ���U  P Some_stuffs_Some_stuffs_ �U  P#��U  $��U  �$��U  �%��U  ��w�.��X /      Workout     P� ��U  �� ��U  �� This_stuffs_This_stuffs_ �U  `� ��U   � ��U  �� ��U  �� ��U  @</�ݡ.(�Y /       Birthday    �� ��U  � ��U  Ы This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `� ��U  �|����.;�Y /      Some_stuffs �'��U   (��U  �(justforfun_justforfun_ ��U  �+��U  �,��U   -��U  �-��U  A��+�.��Y /       Birthday    ����U  p���U  ��This_stuffs_This_stuffs_ �U  @���U   ���U  ����U   ���U  q^p|�.�tZ /       Appointment ���U   ��U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  A�E��.�kg /      Workout     o��U  �o��U  �~Some_stuffs_Some_stuffs_ �U  `r��U   s��U  �s��U  `t��U  �ZR�(�.D�g /       Meeting �U  P���U  ���U  ЮThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  Y�ˇ��.�Vh /       Workout     �� ��U  `� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0� ��U  i �D��.�zh /      Birthday    `_ ��U   ` ��U  `d Some_stuffs_Some_stuffs_ �U  �n ��U  Po ��U  �t ��U  �v ��U  1�(߫.��h /       Birthday    ����U  ���U  гThis_stuffs_This_stuffs_ �U  ���U  ж��U  ����U  P���U  �h�p�.`�h /       Birthday     ���U  ����U  `�This_stuffs_This_stuffs_ �U  ����U  ����U  `���U  ����U  i�j�'�.;i /      Workout      ���U  ����U  `�This_stuffs_This_stuffs_ �U   ���U  ����U    ��U  � ��U  ����^�.�ei /      Meeting      G��U  �G��U   HThis_stuffs_This_stuffs_ �U  �I��U  �J��U  `K��U   L��U  ��Yaz�.��i /       Meeting     �� ��U  @� ��U  0� justforfun_justforfun_  ��U  0� ��U  �� ��U  �� ��U  P� ��U  q1�⭬.3�i /       Appointment ���U  ����U  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �N�=�.�Nu /       Some_stuffs ���U  б��U  ��justforfun_justforfun_ ��U  ���U  ����U  ���U  ж��U  �o"�õ.��w /       Meeting     ���U   ��U  �This_stuffs_This_stuffs_ �U  `��U   ��U  ���U  ���U  i�~'�.�5x /       Workout     �i��U  `j��U   kSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   p��U  pJ�s�.��x /       Workout     � ��U  � ��U  � justforfun_justforfun_  ��U   ! ��U  �! ��U  P% ��U  & ��U  Y;W��.�oy /      Meeting                        Some_stuffs_Some_stuffs_                                     �xb�*�.�y /      Workout     ����U  @���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  A\*��.Pz� /       Workout                        This_stuffs_This_stuffs_                                     YNS�Y�.�� /       Workout     �i��U  `j��U   kjustforfun_justforfun_ ��U  @n��U  �n��U  @o��U   p��U  �8���.[_� /       Workout     �O��U  pP��U  �Pjustforfun_justforfun_ ��U  pS��U  0T��U  �T��U  0U��U  ]+�ٿ.�׆ /      Workout     ���U  й��U  P�justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  ���U  q���.�"� /       Appointment �
��U   ��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ��U  �F̨)�.`L� /       Appointment �=��U  �>��U  `?This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �C��U  P�G���.j� /       Appointment �7 ��U  �8 ��U  @< justforfun_justforfun_ _ �U  pE ��U  0F ��U   J ��U  �J ��U  ۄ o�.qՓ /       Appointment 0����U  ����U  ���justforfun_justforfun_ ���U   ����U  �����U  �����U  p����U  I�P���.E�� /       Appointment `@��U   A��U  �ASome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  `F��U  ���.��� /      Appointment P���U  ����U  ��This_stuffs_This_stuffs_ �U  ���U  ����U  ����U  P���U  q!X?�.�� /       Birthday    `���U  ����U  `�Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  @���U  X����.�� /       Appointment                    Some_stuffs_Some_stuffs_                                     B�P�.�ŗ /      Birthday U  �� ��U  `� ��U   � This_stuffs_This_stuffs_ �U  0� ��U  � ��U  p� ��U  0� ��U  a1x�]�.;B� /       Workout �U  ����U  ���U  Юjustforfun_justforfun_ ��U  ����U  @���U  ���U  ����U  �6h���.j_� /       Workout     ����U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �9��.�ң /       Appointment `w��U  �w��U  �xSome_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  `}��U  ��;y?�.%� /       Meeting     P% ��U  & ��U  �) justforfun_justforfun_  ��U  P3 ��U  4 ��U  �7 ��U  �8 ��U  a��W�.>L� /       Some_stuffs �����U  �����U  ���justforfun_justforfun_ ���U  �����U  @����U  �����U  @����U  p��B��. /       Workout     �� ��U  p� ��U  0� This_stuffs_This_stuffs_ �U   � ��U  �� ��U  �� ��U  @� ��U  s� ��.� /       Workout     ����U  @���U   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ����.�� /      Workout �U  �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U  #���.�:� /      Birthday    ���U   ���U  ��Some_stuffs_Some_stuffs_ �U  `���U   ���U  ����U  ����U  1W�@&�.��� /       Some_stuffs �� ��U  @� ��U  `� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   � ��U  QP��s�.�� /       Birthday nt �?��U  0@��U  �@This_stuffs_This_stuffs_ �U  �B��U  0C��U  �C��U  0D��U  A�.���.N� /       Some_stuffs 0���U  ����U  0�Some_stuffs_Some_stuffs_ �U  0���U  ����U  p���U  ���U  x�3�.� /      Meeting     �� ��U  P� ��U   � This_stuffs_This_stuffs_ �U  0� ��U  � ��U  �� ��U  p� ��U  i��CV�.�h� /      Some_stuffs �I��U  �J��U  `Kjustforfun_justforfun_ ��U   N��U  �N��U  `O��U  �O��U  �Fͪ��.�� /       Birthday U   x��U  �x��U  �yThis_stuffs_This_stuffs_ �U   |��U  �|��U  �}��U  @~��U  �����.�-� /       Appointment � ��U  Ж ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @� ��U  !�7���.�P� /       Birthday    �t��U  �u��U   vThis_stuffs_This_stuffs_ �U  �x��U  `y��U  �y��U  �z��U  �#+�.�t� /       Workout     f��U  �f��U  Pgjustforfun_justforfun_ ��U  j��U  �j��U  �k��U  l��U  �*�#�.��� /      Meeting �U  ����U  @���U   �Some_stuffs_Some_stuffs_ �U  ����U  @���U  ����U  @���U  0��>�.�Ǵ /       Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             ���`U�.�� /       Some_stuffs ���U  `��U   This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @#��U  ��W��.N�� /       Workout     �� ��U  P� ��U   � This_stuffs_This_stuffs_ �U  �� ��U  �� ��U  � ��U  `� ��U  ������.}�� /       Birthday                       This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_             !n����.�۵ /      Meeting �U  ����U   ���U   �Some_stuffs_Some_stuffs_ �U  `���U   ���U  ����U  ����U  �&X�.q� /      Appointment �<��U  p=��U  �=This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �A��U  ��W��.^ƶ /       Birthday nt �� ��U  � ��U  Ы Some_stuffs_Some_stuffs_ �U   � ��U  � ��U  �� ��U  `� ��U  I�l_2Q2 &/      Some_stuffs  ���U  ����U  `�justforfun_justforfun_ ��U  ����U  @���U  ����U  p���U   &��3_2d_ &/       Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             i"�u�_2Sr&/       Workout �U   o��U  �o��U   pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Pt��U  �4`2�&/       Meeting      5��U  �5��U  �6Some_stuffs_Some_stuffs_ �U  `9��U  �9��U  �:��U  `;��U  �]��`2+�&/       Birthday    ����U   ���U  ��justforfun_justforfun_ _ �U  ����U   ���U  ����U   ���U  �}PN`2f&/       Appointment  ���U  ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ���Sa2�&/       Appointment  ��U  ���U  @This_stuffs_This_stuffs_ �U  @��U   ��U  ���U  ���U  H�̙a2�F&/      Meeting     �� ��U  �� ��U   � Some_stuffs_Some_stuffs_ �U  �� ��U  �� ��U  @� ��U   � ��U   �7rbi2��&/      Appointment ���U  `��U   justforfun_justforfun_ ��U  �
��U  ���U  �"��U  @#��U  `U��i2�<&/      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��&��i2>e&/       Workout     ���U  ����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  9�u�i2��&/       Birthday    �t ��U  �v ��U  �z Some_stuffs_Some_stuffs_ �U  �� ��U  P� ��U   � ��U  �� ��U  y0\j2��&/       Birthday    �.��U  `/��U   0This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �4��U  :I��j2{�&/       Birthday fs �$��U  �%��U  P&This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U   +��U  ��v�j2n�&/       Workout     �m��U  `n��U   oSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   s��U  a�E�j2e�&/       Workout     ���U  ���U  pSome_stuffs_Some_stuffs_ �U  p��U  ���U  ���U  p��U  ١���j2�&/       Appointment  J ��U  �J ��U  �N Some_stuffs_Some_stuffs_ �U  �Z ��U  p[ ��U  `_ ��U   ` ��U  i+6k2Ҋ&/       Workout     Ю��U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  ���kk2�&/       Workout �U  �z ��U  �{ ��U  0� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @� ��U  5l!�k2A�&/      Appointment �����U  �����U  ���justforfun_justforfun_ ���U  �����U  @����U  �����U  @����U  yo�s2n&/       Appointment ����U  ����U  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��¯s2U&/       Appointment `� ��U   � ��U  �� Some_stuffs_Some_stuffs_ �U  �� ��U  �� ��U  �� ��U  �� ��U  ��@dt2��&/       Appointment �� ��U  @� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P� ��U  aI�X�t2T� &/       Some_stuffs �_��U  �`��U   ajustforfun_justforfun_ ��U  �c��U  `d��U  �d��U  `e��U  i!Lնt2�� &/       Workout     �� ��U  @� ��U  `� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `� ��U  @U�v�t2!&/      Meeting                        Some_stuffs_Some_stuffs_                                     ْ�+�t2�(!&/       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             A ���u2d9"&/       Meeting     ���U   ��U  �justforfun_justforfun_ ��U  �B��U  pC��U  ` ��U  � ��U  �kF�v2[�"&/       Birthday    ���U  ���U  @Some_stuffs_Some_stuffs_ �U  ���U  0��U  ���U  `	��U  �ةc}20�-&/      Appointment �����U  `����U  ��Some_stuffs_Some_stuffs_ �U  �����U  p����U  0����U  ����U  �}7p�}2�H.&/      Birthday    0� ��U  �� ��U  �� This_stuffs_This_stuffs_ �U  �� ��U  p� ��U  0� ��U   � ��U  �����}2��.&/      Meeting �U  �� ��U  p� ��U  0� justforfun_justforfun_  ��U   � ��U  �� ��U  �� ��U  @� ��U  ���l�}2�.&/      Birthday    �� ��U  P� ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @� ��U  99ck2��0&/      Birthday    p���U  P���U  �justforfun_justforfun_ ��U  Б��U  P���U  В��U  ����U  �q�X�2}1&/       Some_stuffs  ��U  ���U   justforfun_justforfun_ ��U  ���U  @��U   ��U  ���U  �h�2?�1&/      Appointment `��U   ��U  �This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  ���U   ��,4�2�?2&/       Birthday    0����U  ����U  ���Some_stuffs_Some_stuffs_ �U   ����U  �����U  �����U  p����U  0��RN�2&g2&/       Some_stuffs   ��U  � ��U   ! This_stuffs_This_stuffs_ �U  �) ��U  P* ��U  �. ��U  �/ ��U  �T��2?�=&/      Some_stuffs Б��U  P���U  ВSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  �X��d�2�>&/       Birthday U  ����U   ���U  ��justforfun_justforfun_ ��U  ���U   ��U  ����U   ���U  ��n��2~?&/       Some_stuffs �����U  �����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  �&�;Ɉ2??&/      Meeting     �3��U  �4��U   5This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @9��U  y����2ne?&/       Meeting     ����U  0���U  ��justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  p���U  Y8,���2+�?&/       Appointment `O��U  �O��U  �PSome_stuffs_Some_stuffs_ �U  `S��U   T��U  �T��U  Pc��U  i���O�2��?&/       Workout     �7 ��U  �8 ��U  @< Some_stuffs_Some_stuffs_ �U  pE ��U  0F ��U   J ��U  �J ��U  InUc��2Fv@&/       Appointment �����U  `����U  ��Some_stuffs_Some_stuffs_ �U  �����U  p����U  0����U  ����U   }`3�2�ZA&/       Meeting     ���U  ���U  @This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `	��U  �No�L�2ځA&/       Birthday U  ���U  0��U  �Some_stuffs_Some_stuffs_ �U  `��U   ��U  ���U  `��U  �Ew4f�2�A&/       Some_stuffs  J ��U  �J ��U  �N This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ` ��U  y�2�}L&/       Workout     �����U  @����U  ���Some_stuffs_Some_stuffs_ �U  �����U  P����U  �����U  @����U  p�����2N!M&/       Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             )z��-�2�kM&/       Appointment  j��U  �j��U  `kSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �o��U  �'ٙ�2��O&/       Birthday U  Б��U  P���U  ВThis_stuffs_This_stuffs_ �U  P���U  ���U  ����U  P���U  �*�4�2�yP&/       Some_stuffs P���U  ���U  лThis_stuffs_This_stuffs_ �U  P���U  ���U  ����U  ���U  q���j�2U�P&/      Appointment  ���U  ����U  @�Some_stuffs_Some_stuffs_ �U  ����U  ����U   ���U  ����U  ���S-�2�\&/       Birthday    �� ��U  �� ��U  P� justforfun_justforfun_  ��U  �� ��U  @� ��U  `� ��U   � ��U  ��c~�2@�\&/       Workout     @���U  ����U  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  !K���2��]&/       Workout ffs � ��U  ���U  Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �x |�2��^&/       Appointment Ѕ��U  ����U  @�This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  h��Ŵ�2�^&/      Birthday                       Some_stuffs_Some_stuffs_                                     ��0;�2,l_&/       Workout     �� ��U  @� ��U  �� This_stuffs_This_stuffs_ �U  � ��U  Щ ��U  �� ��U  � ��U  H6ށ�2	`&/      Birthday    p� ��U  �� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   � ��U   �v��2�Qk&/       Meeting     � ��U  � ��U  � Some_stuffs_Some_stuffs_ �U   ! ��U  �! ��U  P% ��U  & ��U  ��tz{�28l&/       Birthday    л��U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  i�H�G�2�Pm&/       Some_stuffs                    Some_stuffs_Some_stuffs_                                     A&eHz�2~�m&/       Meeting     ���U  ����U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  (l벧2��m&/       Workout     м ��U  �� ��U  P� justforfun_justforfun_  ��U  P� ��U  � ��U  �� ��U  �� ��U  YK��2�6n&/      Birthday nt �����U  �����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  8����2�n&/       Birthday    P����U  ����U  P��Some_stuffs_Some_stuffs_ �U  P����U  ����U  �����U  @����U  y�K�f�2so&/      Some_stuffs ���U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ���+�2Z�z&/       Workout     �|��U  `}��U  ��This_stuffs_This_stuffs_ �U  ����U  `���U   ���U  ����U  QL�F^�2	{&/       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �s<��2b�{&/       Some_stuffs �3��U  �4��U   5This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @9��U  �X�F�2~ |&/      Meeting                        justforfun_justforfun_                                       �v�a�2��|&/       Birthday    ����U  @���U   �This_stuffs_This_stuffs_ �U  ����U  ����U  @���U   ���U  aV줯�2y	}&/       Birthday    p���U  0���U  ��justforfun_justforfun_ ��U  ����U  ����U  p���U  P���U  s�d0�2��}&/      Workout �U  �����U  �����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  ���.Ͳ2��~&/       Birthday nt �4��U  �5��U  p6justforfun_justforfun_ _ �U  �8��U  p9��U  �9��U  p:��U   �V�)�2D؉&/       Some_stuffs `H��U   I��U  �Ijustforfun_justforfun_ _ �U  �L��U  `M��U  �M��U  �N��U  ��&�_�2Z*�&/       Workout     ���U  ����U  �This_stuffs_This_stuffs_ �U  ���U  й��U  P���U  ���U  )q+��2��&/      Some_stuffs  v��U  �v��U  `wjustforfun_justforfun_ ��U  �y��U  �z��U  `{��U  �{��U  �q���2S=�&/       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_             ��PI�2g��&/      Meeting     ����U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p���U  vs���28��&/      Some_stuffs �� ��U  p� ��U  0� justforfun_justforfun_  ��U   � ��U  �� ��U  �� ��U  @� ��U  ���s�2�[�&/       Birthday    ����U  ����U   �justforfun_justforfun_ ��U  ����U  ����U  ����U  @���U  (X:��2E��&/       Workout     � ��U  � ��U  � justforfun_justforfun_  ��U   ! ��U  �! ��U  P% ��U  & ��U  �:*��2���&/       Some_stuffs  � ��U  �� ��U  @� justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  �� ��U  pHA��2�ј&/      Appointment �����U  `����U  ��This_stuffs_This_stuffs_ �U  �����U  p����U  0����U  ����U  ��⫧�2h��&/       Meeting     ���U  И��U  ��This_stuffs_This_stuffs_ �U  ����U  ���U  Ю��U  P���U  ѽ���2Cۙ&/       Appointment �S ��U  �U ��U  �Z This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0j ��U  g���2S�&/       Workout     �7 ��U  �8 ��U  @< Some_stuffs_Some_stuffs_ �U  pE ��U  0F ��U   J ��U  �J ��U  )�����2�f�&/       Workout     ����U   ���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  AU����2g��&/       Workout     e��U  �e��U  fThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �j��U  8�YA1�2'�&/      Workout     P���U  ���U  ��This_stuffs_This_stuffs_ �U  ����U   ���U  ����U  @���U  0`�E�2f%�&/       Meeting                        justforfun_justforfun_                                       �����2\��&/       Birthday    �:��U  `;��U   <Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �A��U  �z����2��&/       Some_stuffs �Z��U   [��U  �[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �`��U  ����2��&/       Some_stuffs Ы ��U  �� ��U  P� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  � ��U  )C4��2<�&/       Some_stuffs �7 ��U  �8 ��U  @< justforfun_justforfun_  ��U  pE ��U  0F ��U   J ��U  �J ��U  Y�-�&�2E�&/       Meeting     `� ��U   � ��U  �� This_stuffs_This_stuffs_ �U  �� ��U  �� ��U  �� ��U  �� ��U  9�]A�2H;�&/       Birthday nt 0b��U  �b��U  �cThis_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  h��U  ��a��2ԧ�&/       Workout �U  ����U  `���U  �This_stuffs_This_stuffs_ �U  ���U  б��U  ����U  ���U  `R7/��2l��&/       Appointment �����U  �����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @����U  �Йn-�2{��&/      Workout                        Some_stuffs_Some_stuffs_                                     *��\�2��&/       Meeting �U  �P��U  `Q��U   Rjustforfun_justforfun_ ��U  �T��U  Pc��U  �V��U  �W��U  @����2~�&/       Workout                        justforfun_justforfun_                                       ɱ�!��2Ҫ&/       Some_stuffs ����U  @���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  qǬk`�26i�&/       Appointment �� ��U  �� ��U  � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  `�PJ��2̵�&/       Birthday    �� ��U  `� ��U   � This_stuffs_This_stuffs_ �U  0� ��U  � ��U  p� ��U  0� ��U  ��u��2��&/      Appointment 0����U  ����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p����U  ������,��/       Some_stuffs �� ��U  @� ��U  `� justforfun_justforfun_  ��U  �� ��U  �� ��U  `� ��U   � ��U  ������,�/       Meeting      5��U  �5��U   6This_stuffs_This_stuffs_ �U  �8��U  @9��U  `R��U   S��U  !%�3�F�,�$/       Meeting     `���U  ����U  ��justforfun_justforfun_ ��U  ����U  `���U  ����U  ����U  "%�3�F�,�$/      Some_stuffs ���U  p���U  �This_stuffs_This_stuffs_ �U  0���U  ���U  ����U  p���U  �O�?Qn�,f9%/       Workout     0����U  ����U  ���Some_stuffs_Some_stuffs_ �U   ����U  �����U  �����U  p����U  �O�?Qn�,A%/       Some_stuffs �|��U  `}��U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ���B;�,�'/      Workout �U  ����U  @���U  ��This_stuffs_This_stuffs_ �U   ���U  ����U  @���U   ���U  ���B;�,�'/       Meeting ent @7��U   8��U  �8This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U   =��U  ��]�,�3/       Birthday    `O��U  �O��U  `PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �U��U  ��]�,�$3/      Meeting     �����U  @����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @����U  �C�bu-�,��3/       Workout     0%��U  �%��U  p&justforfun_justforfun_ ��U  �(��U  p)��U  �)��U  p*��U  A��l�T�,�U4/       Meeting     ���U   ��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @��U  B��l�T�,xY4/       Workout     p{��U  �{��U  p|This_stuffs_This_stuffs_ �U   ��U  ���U  P���U  Ѐ��U  ����,�|6/      Birthday     A��U  �A��U  �BThis_stuffs_This_stuffs_ �U  �E��U  `F��U   G��U  �G��U  ����,$|6/       Appointment `���U  ���U  ��justforfun_justforfun_ ��U  ���U  ����U  ���U  б��U  `c�%[*�,l*C/       Appointment м ��U  �� ��U  P� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  y"A涥,�GE/      Appointment �� ��U  � ��U  Ы justforfun_justforfun_  ��U   � ��U  � ��U  �� ��U  `� ��U  z"A涥,�FE/       Meeting     �� ��U  @� ��U  `� justforfun_justforfun_  ��U  �� ��U  �� ��U  `� ��U   � ��U  !����ե,��E/       Meeting     P���U  ���U  ��This_stuffs_This_stuffs_ �U  ��U  ���U  @��U  ���U  "����ե,��E/       Workout     ���U  ����U  �justforfun_justforfun_ ��U  P���U  ����U  ����U  ���U  ��?�ߥ,��E/       Some_stuffs P� ��U  p� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  ��?�ߥ,&�E/       Some_stuffs 0� ��U  � ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  �#p���,�[F/      Some_stuffs �����U  �����U  ���Some_stuffs_Some_stuffs_ �U  �����U  @����U  �����U  @����U  �#p���,YF/       Meeting     �d��U  `e��U  �eThis_stuffs_This_stuffs_ �U  `h��U   i��U  �i��U  `j��U  If"k��,��Q/       Birthday fs �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U  Jf"k��,~�Q/      Meeting                        justforfun_justforfun_                                       Q|4�b�,xS/       Birthday    0����U  ����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p����U  R|4�b�,�vS/       Some_stuffs P���U  ����U  ��justforfun_justforfun_ ��U   ���U  ����U  ����U  @���U  ���x_l�,��S/       Birthday U  �����U  �����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  i���,�9a/       Birthday                       Some_stuffs_Some_stuffs_                                     j���,:5a/       Some_stuffs ����U  P���U  �justforfun_justforfun_ ��U  ����U  ����U  P���U  ����U  �4p{R�,'�b/       Some_stuffs ����U  ���U  ЮThis_stuffs_This_stuffs_ �U  ����U  @���U  ���U  ����U  �4p{R�,վb/      Some_stuffs `��U  ���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `��U  i顸Q]�,t�b/       Workout     0b��U  �b��U  �cSome_stuffs_Some_stuffs_ �U  f��U  �f��U  Pg��U  h��U  j顸Q]�,��b/       Appointment ���U   ��U  �justforfun_justforfun_ _ �U  �B��U  pC��U  ` ��U  � ��U  Q8V��f�,�
c/       Appointment �� ��U  p� ��U  0� Some_stuffs_Some_stuffs_ �U   � ��U  �� ��U  �� ��U  @� ��U  R8V��f�,5c/       Appointment 0����U  ����U  ���This_stuffs_This_stuffs_ �U   ����U  �����U  �����U  p����U  Av�Q�˰,�-p/      Appointment � ��U  Ж ��U  �� This_stuffs_This_stuffs_ �U   � ��U  �� ��U  �� ��U  @� ��U  Bv�Q�˰,�-p/       Meeting     �(��U  p)��U  �)This_stuffs_This_stuffs_ �U  0,��U  �,��U  p-��U  0.��U  �5���,�=q/      Some_stuffs 0����U  ����U  ���This_stuffs_This_stuffs_ �U   ����U  �����U  �����U  p����U  I����9�,��q/      Appointment                    justforfun_justforfun_                                       J����9�,b�q/       Workout     �t ��U  �v ��U  �z This_stuffs_This_stuffs_ �U  �� ��U  P� ��U   � ��U  �� ��U  )D8Xm�,&�r/       Meeting �U  �����U  �����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @����U  *D8Xm�,��r/      Workout     �����U  ����U  ���justforfun_justforfun_  ��U  � ��U  @	 ��U  P ��U   ��U  ��+ѱ,]t/       Workout     �]��U  p^��U  0_Some_stuffs_Some_stuffs_ �U  0b��U  �b��U  �c��U  Pd��U  i2�4ݱ,�Jt/       Some_stuffs  ���U  ����U  @�Some_stuffs_Some_stuffs_ �U  ����U  ����U  @���U   ���U  j2�4ݱ,�Dt/      Some_stuffs ����U  P���U  �Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  П��U  Q��J2ƴ,��/       Meeting ffs p\��U  0]��U  �]This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �b��U  R��J2ƴ,�/      Some_stuffs  6��U  �6��U  @7justforfun_justforfun_ ��U  `R��U   S��U   ;��U  �;��U  q�F�l�,�-�/       Workout     �� ��U  `� ��U   � Some_stuffs_Some_stuffs_ �U  0� ��U  � ��U  p� ��U  0� ��U  r�F�l�,.�/       Appointment `��U  ���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @��U  �l�|�,���/       Birthday    `R��U   S��U   ;Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �?��U  �l�|�,Ȩ�/      Meeting     �� ��U  p� ��U  0� This_stuffs_This_stuffs_ �U  @� ��U   � ��U  �� ��U  �� ��U  �� ���,�ˀ/       Workout �U  ����U  ����U  P�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �� ���,�ˀ/       Birthday U  `���U   ���U  ��justforfun_justforfun_ ��U    ��U  � ��U  `��U  ���U  �~4��!�,���/       Appointment �� ��U  � ��U  Ы Some_stuffs_Some_stuffs_ �U   � ��U  � ��U  �� ��U  `� ��U  X7�O�@�,�g�/      Meeting �U  �� ��U  p� ��U  0� Some_stuffs_Some_stuffs_ �U   � ��U  �� ��U  �� ��U  @� ��U  Гw�͵,���/       Meeting     �����U  p����U  0��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �����U  Q��]q��,�׎/       Meeting     �� ��U  `� ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  R��]q��,֎/       Workout     0-��U  �-��U  p.This_stuffs_This_stuffs_ �U  �0��U  �1��U  02��U  �2��U  A�<�,?o�/       Some_stuffs �����U  �����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  B�<�,�r�/      Appointment �"��U  @#��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U   !P�[�,�J�/       Some_stuffs                    Some_stuffs_Some_stuffs_                                     !��_�o�,3��/      Birthday    `��U   ��U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �:��U  "��_�o�, ��/       Birthday    P���U  Ё��U  P�This_stuffs_This_stuffs_ �U  ����U  ���U  Ѕ��U  ����U  �.�K��,�Z�/       Appointment �����U  @����U  ���Some_stuffs_Some_stuffs_ �U  �����U  P����U  �����U  @����U  !��ե��,�e�/      Meeting     �N��U  pO��U  �OThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0T��U  "��ե��,Ih�/       Appointment �E��U  `F��U   GThis_stuffs_This_stuffs_ �U  �U��U  pV��U  �I��U  �J��U  9\���U�,ʱ�/       Some_stuffs  H��U  �H��U  �USome_stuffs_Some_stuffs_ �U  `K��U   L��U  �L��U  `M��U  :\���U�,歠/      Some_stuffs ���U  ����U  оSome_stuffs_Some_stuffs_ �U  ���U  ����U  @���U  ����U  qöќ��,8n�/       Workout     �� ��U  p� ��U  �� justforfun_justforfun_ _Some_stuffs_Some_stuffs_ �U  �� ��U  röќ��,qr�/       Meeting     @���U  ����U  ��This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  @���U  �y�	z�,v��/      Birthday    P% ��U  & ��U  �) Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �8 ��U  �y�	z�,���/       Some_stuffs ���U  P��U   Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `"��U  Y)Ġ��,�/      Some_stuffs  g��U  �g��U  `hSome_stuffs_Some_stuffs_ �U   k��U  �k��U   m��U  �m��U  Z)Ġ��,`��/       Appointment p� ��U  0� ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  �Ȩ���,�w�/      Workout     ����U  @���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  �Ȩ���,lu�/       Workout �U  ����U  @���U  ��Some_stuffs_Some_stuffs_ �U  ����U   ���U  ����U  ����U  �����,��/       Appointment ����U  P���U  ��justforfun_justforfun_ ��U  ����U   ���U  ����U  `���U  �����,�/      Meeting     � ��U  � ��U  � This_stuffs_This_stuffs_ �U  0 ��U  � ��U  � ��U  � ��U  ��T�0��,0��/       Some_stuffs ���U  ���U  P Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �%��U  q���-�9� /       Birthday    �l��U  Pm��U  �mThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �q��U  r���-i<� /      Meeting ffs �����U  `����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  s���-=8� /       Appointment  |��U  �|��U  �}This_stuffs_This_stuffs_ �U  @���U  ����U  @���U   ���U  t���-8� /       Some_stuffs ����U  ����U   �Some_stuffs_Some_stuffs_ �U  ����U  `���U   ���U  ����U  �	{J�#.8
 /       Meeting     �����U  p����U  p��Some_stuffs_Some_stuffs_ �U  @����U  ����U  P����U  ����U  �	{J�#.:y
 /      Workout     �� ��U  P� ��U  �� justforfun_justforfun_  ��U  �� ��U  �� ��U   � ��U  �� ��U  ����̏#."�
 /       Some_stuffs �Y��U  �Z��U  0[This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  �_��U  ����̏#.֟
 /       Birthday fs �G��U  0H��U  �HThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �L��U  ����#.j /       Meeting �U  ����U  @���U   �Some_stuffs_Some_stuffs_ �U  ����U   ���U  ����U  ����U  ����#.[ /       Appointment p/��U  00��U  �0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �5��U  !���#.�� /      Workout     �� ��U  p� ��U  0� justforfun_justforfun_  ��U   � ��U  �� ��U  �� ��U  @� ��U  "���#.5� /       Birthday    `���U  ����U  ��Some_stuffs_Some_stuffs_ �U  ����U   ���U  ����U  ����U  q��:$.�9 /       Some_stuffs ����U   ���U  ��Some_stuffs_Some_stuffs_ �U  ����U  ����U   ���U  ����U  r��:$.e= /       Birthday    ����U  `���U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  ͂��Y$.� /       Workout �U  ���U  0��U  �justforfun_justforfun_ ��U  `��U   ��U  ���U  `��U  ͂��Y$.� /      Appointment �����U  @����U   ��Some_stuffs_Some_stuffs_ �U  �����U  �  ��U  � ��U  � ��U  �#���b$.�� /       Appointment �����U  �����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  q�y���$.�N /      Some_stuffs �T��U  Pc��U  �VThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �[��U  r�y���$.FM /       Workout     `?��U  �?��U  `@Some_stuffs_Some_stuffs_ �U   C��U  �C��U  `D��U  �D��U  ��)\3�$.4� /       Meeting     ����U  @���U  ��Some_stuffs_Some_stuffs_ �U  ����U  @���U  ����U  @���U  ٷ:��'.�� /       Some_stuffs ���U  `��U   This_stuffs_This_stuffs_ �U  ���U  `��U  ���U  ���U  ڷ:��'.�� /       Some_stuffs ���U  `���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �_= �'.�� /       Meeting      $��U  �$��U   %This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P)��U  �_= �'.� /       Birthday    ���U  ���U  P Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �%��U  ��"�O�'.w� /      Appointment �+��U  �,��U   -This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �=��U   IE���'.�G /       Some_stuffs ����U  ����U  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  ����(.l, /      Workout �U  �
��U  ���U  �"justforfun_justforfun_ ��U   ��U  ���U   ��U  ���U  ����(.2 /       Birthday     ��U  ���U   Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @��U  9��sA(.'� /       Workout     �� ��U  p� ��U  0� Some_stuffs_Some_stuffs_ �U  0� ��U   � ��U  �� ��U  �� ��U  :��sA(.s� /       Some_stuffs `K��U   L��U  �LSome_stuffs_Some_stuffs_ �U  `O��U  �O��U  `P��U   Q��U  x�H��J(.� /       Workout �U    ��U  � ��U  `!Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �%��U  	a�T(.� /       Meeting      5��U  �5��U   6Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   S��U  
a�T(._ /       Meeting �U  P���U  У��U  ��Some_stuffs_Some_stuffs_ �U  ����U  @���U  ����U  ����U  �uo�Qr(.h� /       Workout �U  �t��U  �u��U   vSome_stuffs_Some_stuffs_ �U   x��U  �x��U  �y��U  @z��U  �uo�Qr(.�� /       Workout �U  @���U   ���U  ��justforfun_justforfun_ ��U  p���U  ���U  ����U   ���U  ��2s�+.��) /       Workout     ����U  ����U  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ��2s�+.��) /       Some_stuffs  %��U  �%��U   &This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P*��U  �OgP/.�8 /       Workout     ����U  p���U  ��This_stuffs_This_stuffs_ �U  @���U   ���U  ����U   ���U  �OgP/.�8 /       Birthday fs @��U  ���U  @justforfun_justforfun_ _ ome_stuffs_Some_stuffs_ �U  ���U  1�kt�m/.C�8 /      Some_stuffs  C��U  �C��U  `DSome_stuffs_Some_stuffs_ �U  �F��U  �G��U  `H��U   I��U  2�kt�m/.��8 /       Workout      � ��U  �� ��U  �� justforfun_justforfun_  ��U   � ��U  �� ��U  �� ��U  @� ��U  a�6-0.�u; /       Workout     �����U  @����U   ��This_stuffs_This_stuffs_ �U  �����U  �  ��U  � ��U  � ��U  b�6-0.w; /       Workout     ���U  0��U  �Some_stuffs_Some_stuffs_ �U  `��U   ��U  ���U  `��U  ��]#&L3.G�G /       Meeting     `*��U   +��U  �+This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �0��U  ��]#&L3..�G /      Birthday    p&��U  �&��U  �'This_stuffs_This_stuffs_ �U  �)��U  p*��U  �*��U  p+��U  hM�G1�3.M�H /       Some_stuffs �~��U   ��U  �pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �u��U  �]+�ٯ3.�I /       Meeting     ���U  ����U  p�Some_stuffs_Some_stuffs_ �U  p���U  0���U  ����U  ����U  �]+�ٯ3.�I /       Birthday    `9��U  �9��U  �:justforfun_justforfun_ ��U  `>��U  �>��U  �?��U  `@��U  (^~2�3.��I /       Birthday U  ���U  ���U  pThis_stuffs_This_stuffs_ �U  p��U  ���U  ���U  p��U  �;�G4.�XK /      Meeting     �� ��U  p� ��U  0� justforfun_justforfun_  ��U   � ��U  �� ��U  �� ��U  @� ��U  �;�G4.CVK /       Appointment �����U  ����U  ���Some_stuffs_Some_stuffs_ �U  � ��U  @	 ��U  P ��U   ��U  ��P[4.͢K /       Birthday    п��U  P���U  �Some_stuffs_Some_stuffs_ �U  ���U  ����U  P���U  ����U  ��P[4.N�K /      Meeting     �� ��U  �� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `� ��U  �*Ү�7.�NX /      Workout ent 0����U  ����U  ���justforfun_justforfun_ ���U   ����U  �����U  �����U  p����U  �*Ү�7.rJX /       Some_stuffs 0-��U  �-��U  p.justforfun_justforfun_ _ his_stuffs_This_stuffs_ �U  �2��U  ��O�7.��X /       Birthday     ���U  ����U  `�Some_stuffs_Some_stuffs_ �U   ���U  ����U    ��U  � ��U  ��O�7.��X /      Workout     �Q��U  �l��U  �SThis_stuffs_This_stuffs_ �U  �V��U  `W��U  �W��U  �X��U  A}+0��7.$�Y /       Workout     ���U   ��U  �Some_stuffs_Some_stuffs_ �U   ��U  ���U   ��U  ���U  B}+0��7.x�Y /       Workout     ����U  ����U  `�justforfun_justforfun_ ��U  ����U   ���U  ����U  `���U  �}Gw$8.cGZ /       Appointment 0� ��U  �� ��U  �� This_stuffs_This_stuffs_ �U  �� ��U  @� ��U  �� ��U  �� ��U  �dl��<.	�i /       Birthday nt ���U  ���U  P Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �%��U  �dl��<.��i /      Appointment ����U  P���U  �Some_stuffs_Some_stuffs_ �U  ���U  Л��U  ����U  ���U  q��CN�?.�x /       Some_stuffs ����U  P���U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  r��CN�?.��x /       Some_stuffs ���U  `���U  �This_stuffs_This_stuffs_ �U  ����U  `���U   ���U  ����U  @��3:@.(�y /      Workout                        justforfun_justforfun_                                       �,�E�D@.�y /       Birthday    P% ��U  & ��U  �) Some_stuffs_Some_stuffs_ �U  P3 ��U  4 ��U  �7 ��U  �8 ��U  �,�E�D@.��y /       Birthday    ����U   ���U   �Some_stuffs_Some_stuffs_ �U  `���U   ���U  ����U  ����U  	���+�C.a؆ /       Workout     ���U   ��U  �This_stuffs_This_stuffs_ �U  `��U  ���U  ���U  `��U  
���+�C.�چ /       Workout     �k��U  l��U  �lThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ��U  Q�����C.�� /       Appointment �)��U  �*��U  p+Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p/��U  R�����C.�� /      Some_stuffs ���U  ж��U  ��Some_stuffs_Some_stuffs_ �U  P���U  ���U  л��U  ����U  `OA;$"D.쫈 /       Meeting     P% ��U  & ��U  �) Some_stuffs_Some_stuffs_ �U  P3 ��U  4 ��U  �7 ��U  �8 ��U  Y	_E H.��� /       Appointment ����U  @���U   �This_stuffs_This_stuffs_ �U  ����U   ���U  ����U  ����U  Z	_E H.#�� /       Some_stuffs 0 ��U  � ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �! ��U  ���J	H.�ŗ /       Birthday    0����U  ����U  ���Some_stuffs_Some_stuffs_ �U   ����U  �����U  �����U  p����U  ���J	H.Ǘ /       Appointment В��U  ����U  �This_stuffs_This_stuffs_ �U  ����U  P���U  ���U  И��U  ��i�cK.4�� /       Some_stuffs �� ��U  `� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0� ��U  �=r�&K.\ۣ /       Birthday     ���U  ����U   �This_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  @���U  �=r�&K.�ӣ /      Birthday    0b��U  �b��U  �cSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  h��U  �I�O&1K.4�� /       Some_stuffs �����U  ����U  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ��U  q���ycK.߽� /      Birthday    �����U  `����U  ��This_stuffs_This_stuffs_ �U  �����U  p����U  0����U  ����U  r���ycK.�� /       Some_stuffs ����U  `���U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  y-���O.�� /       Birthday U  �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U  z-���O.�� /       Some_stuffs �����U  p����U  0��Some_stuffs_Some_stuffs_ �U  P����U   ����U   ����U  �����U  ���,�`O.�.� /       Birthday    ���U  ����U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  ���,�`O.�*� /      Appointment ����U  p���U  ��Some_stuffs_Some_stuffs_ �U  p���U  0���U  ����U  0���U  1�%ձ�O.CŴ /       Some_stuffs                    Some_stuffs_Some_stuffs_                                     2�%ձ�O.J˴ /      Some_stuffs �� ��U  @� ��U  `� This_stuffs_This_stuffs_ �U  �� ��U  �� ��U  `� ��U   � ��U  ᔸ�q�O.�� /       Some_stuffs �����U  p����U  p��Some_stuffs_Some_stuffs_ �U  @����U  ����U  P����U  ����U  ┸�q�O.�� /       Meeting     �U��U  pV��U  �ISome_stuffs_Some_stuffs_ �U  �L��U  `M��U   N��U  �N��U  �a��P.]�� /       Meeting ent �� ��U  @� ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  � ��U  Ѽ6���X/��+ /       Meeting  fs �����U  @����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  Ҽ6���X/ȗ+ /       Some_stuffs `!��U  �!��U   :justforfun_justforfun_ ��U  0%��U  �%��U  p&��U  �&��U  Ӽ6���X/}�+ /      Birthday                       justforfun_justforfun_                                       Լ6���X/>�+ /       Some_stuffs �Q��U  �R��U  pSSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pW��U  ռ6���X/��+ /       Appointment �:��U  `;��U   <Some_stuffs_Some_stuffs_ �U  �?��U  `@��U   A��U  �A��U  !��g�/�b &/       Some_stuffs pX��U  0Y��U  �YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  p^��U  "��g�/�\ &/      Workout     ���U  ���U  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p��U  I�ΐ���/6G&/       Workout     ����U  ����U  �This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  J�ΐ���/	@&/       Workout     �. ��U  �/ ��U  P3 justforfun_justforfun_  ��U  @< ��U   = ��U  �@ ��U  �A ��U  �&~|ڮ/�&/       Birthday     � ��U  �� ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  P� ��U  !BK��/,�&/       Some_stuffs P� ��U  @� ��U  0� justforfun_justforfun_ _ �U  0� ��U  �� ��U  �� ��U  p� ��U  "BK��/�&/       Workout     P���U  Ѐ��U  P�This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  ���U  aY.��/s;&/       Birthday                       Some_stuffs_Some_stuffs_                                     bY.��/�:&/       Appointment  ��U  ���U  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @���U  �^�Y��/��&/      Some_stuffs p9��U  0:��U  �:justforfun_justforfun_ ��U  �<��U  p=��U  �=��U  p>��U  �^�Y��/�&/       Birthday    ����U  @���U  ��justforfun_justforfun_ ��U  @���U  ����U  ����U  @���U  	����/L�&/       Birthday    � ��U  � ��U  � This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  & ��U  
����/o�&/       Meeting ffs `���U  ����U  `�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ���U  A�4Y�X�/a!&/       Meeting                        Some_stuffs_Some_stuffs_                                     B�4Y�X�/'!&/       Birthday U  ����U   ���U  �Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  `���U  �F�6ܹ/��.&/       Birthday    @��U   ��U  �justforfun_justforfun_ ��U  ���U  ���U  ���U  0��U  �F�6ܹ/��.&/       Meeting     � ��U  � ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  & ��U  uּ�̺/�@2&/      Appointment pi ��U  0j ��U  �n Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  uּ�̺/eB2&/       Appointment P����U  ����U  P��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @����U  1�y�ֺ/*g2&/       Birthday     N��U  �N��U  `OSome_stuffs_Some_stuffs_ �U   R��U  �R��U  `S��U   T��U  2�y�ֺ/zi2&/      Birthday    ���U  P��U   Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `"��U  !��P��/�aA&/      Workout      ���U  ����U  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  "��P��/�ZA&/       Appointment �V��U  �W��U  pXThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0]��U  �^�.��/Z�A&/       Appointment ���U  ж��U  ��Some_stuffs_Some_stuffs_ �U  P���U  ���U  л��U  ����U  �^�.��/S�A&/       Meeting     ����U  ����U  �This_stuffs_This_stuffs_ �U  ����U  ����U  p���U  0���U  q`u�;��/M&/      Meeting ffs `_ ��U   ` ��U  `d Some_stuffs_Some_stuffs_ �U  �n ��U  Po ��U  �t ��U  �v ��U  r`u�;��/eM&/       Meeting      0��U  �0��U   =Some_stuffs_Some_stuffs_ �U  �3��U  �4��U   5��U  �5��U  	���/��[&/       Meeting     @< ��U   = ��U  �@ Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �O ��U  i+�7�R�/��^&/       Meeting �U  �����U  @����U  ���This_stuffs_This_stuffs_ �U  �����U  P����U  �����U  @����U  j+�7�R�/��^&/       Appointment ����U   ���U  ��Some_stuffs_Some_stuffs_ �U  ����U  @���U  ����U  ����U  IsR���/(`&/       Birthday    ���U  `���U  �This_stuffs_This_stuffs_ �U   ���U  ����U  `���U  ����U  JsR���/`&/       Birthday    ����U   ���U  ��Some_stuffs_Some_stuffs_ ome_stuffs_Some_stuffs_ �U  ����U  !��1���/nXk&/       Workout     �� ��U  `� ��U   � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0� ��U  "��1���/Qk&/      Birthday U  @r��U   s��U  �sThis_stuffs_This_stuffs_ �U   v��U  �v��U   w��U  �w��U  X�����/Kel&/      Workout �U  �����U  �����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  9hcl�`�/�n&/       Workout     @� ��U   � ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P� ��U  :hcl�`�/��n&/       Workout ffs `*��U   +��U  �+Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �0��U  �����/�|&/       Birthday nt P���U  ���U  ��Some_stuffs_Some_stuffs_ his_stuffs_This_stuffs_ �U  ����U  �����/n|&/       Birthday    p|��U  0}��U  �}This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  Ё��U  �����/H�|&/       Appointment P����U  ����U  P��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  �����/d�|&/       Meeting     `���U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  u��S�/W�}&/       Birthday    � ��U  � ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  & ��U  u��S�/��}&/       Appointment ���U  Л��U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @���U  !�n��p�/�ى&/       Workout     ���U  ����U  @�Some_stuffs_Some_stuffs_ �U  ����U   ���U  ����U  @���U  "�n��p�/�݉&/       Meeting ent  ���U  ����U  @�justforfun_justforfun_ ��U  ����U  @���U   ���U  ����U  )5cFAc�/)��&/      Some_stuffs �� ��U  p� ��U  0� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  *5cFAc�/���&/       Meeting �U  ���U  ���U  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p��U  �	;�l�/���&/       Appointment ����U  `���U  ��Some_stuffs_Some_stuffs_ �U  `���U   ���U  ����U  ����U  �	;�l�/˪�&/       Some_stuffs � ��U  ���U  0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  qUt�kO�/�͘&/       Appointment ����U  @���U   �justforfun_justforfun_ ��U  ����U  @���U  ����U  @���U  rUt�kO�/tИ&/       Appointment В��U  ����U  �justforfun_justforfun_ _ �U  ����U  P���U  ���U  И��U  ��Qfc�/8�&/      Some_stuffs                    This_stuffs_This_stuffs_                                     ��Z}.��/�z�&/       Workout                        This_stuffs_This_stuffs_                                     9��Xl#�/���&/       Meeting     0[��U  �[��U  p\Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  pa��U  :��Xl#�/u�&/       Some_stuffs ���U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  1���+�/�%�&/      Some_stuffs @^��U  �^��U  �_Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  Pc��U  2���+�/G&�&/       Birthday    �����U  `����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �*>"K�/h��&/      Appointment @� ��U   � ��U  �� justforfun_justforfun_  ��U  �� ��U   ��U  �� ��U  @ ��U  �*>"K�/.��&/       Meeting     �� ��U  �� ��U  `� justforfun_justforfun_  ��U   � ��U  �� ��U  �� ��U  �� ��U  �7g�/s��&/      Workout     P3 ��U  4 ��U  �7 justforfun_justforfun_  ��U  �@ ��U  �A ��U  pE ��U  0F ��U  �7g�/%��&/       Appointment �)��U  �*��U  p+justforfun_justforfun_ ��U  p-��U  �-��U  �.��U  p/��U  a�u�}�/`��&/       Workout                        This_stuffs_This_stuffs_                                     b�u�}�/���&/       Workout     �l��U  Pm��U  �mjustforfun_justforfun_ ��U  �~��U   ��U  �p��U  �q��U  ��:��/��&/       Some_stuffs �p��U  �q��U  `rSome_stuffs_Some_stuffs_ �U  �t��U  �u��U   v��U  �v��U  ��:��/+��&/       Workout     P���U  ���U  ��This_stuffs_This_stuffs_ �U  ����U  P���U  ���U  Л��U  ɒ5c��/�&/       Workout     `O��U  �O��U  �PSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  Pc��U  ɒ5c��/5�&/       Meeting �U  `���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  A�:����/7~�&/      Meeting                        justforfun_justforfun_                                       B�:����/8��&/       Some_stuffs @���U  ����U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  a.VT1�/ּ�&/       Workout     �� ��U  �� ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  b.VT1�/���&/       Birthday    �c��U  Pd��U  eThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �i��U  ����E�/��&/       Birthday    P� ��U  @� ��U  0� justforfun_justforfun_  ��U  0� ��U  �� ��U  �� ��U  p� ��U  ����E�/n�&/       Birthday    ���U  ���U    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p$��U  	t�T�nV��{&/       Meeting     �3��U  �4��U   5Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �9��U  
t�T�nV6�{&/       Meeting     �� ��U  p� ��U  0� Some_stuffs_Some_stuffs_ �U   � ��U  �� ��U  �� ��U  @� ��U  t�T�nV�{&/       Workout     `@��U   A��U  �AThis_stuffs_This_stuffs_ his_stuffs_This_stuffs_ �U  `F��U  t�T�nVէ{&/       Workout     ���U  @��U   Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  I�"�XƄYR� /       Meeting �U  � ��U  � ��U  � Some_stuffs_Some_stuffs_ �U  0 ��U  � ��U  � ��U  � ��U  J�"�XƄY�� /       Workout     0����U  ����U  ���This_stuffs_This_stuffs_ �U   ����U  �����U  �����U  p����U  K�"�XƄY9� /      Some_stuffs 0b��U  �b��U  �cSome_stuffs_Some_stuffs_ �U  f��U  �f��U  Pg��U  h��U  L�"�XƄY}� /       Appointment В��U  ����U  �This_stuffs_This_stuffs_ �U  ����U  P���U  ���U  И��U  X�\>�cm�'$/      Some_stuffs ���U  ���U  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p��U  �|g��+nE�1&/       Workout                        This_stuffs_This_stuffs_                                     �|g��+n��1&/       Workout �U  �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U  �|g��+n��1&/       Workout     �����U  @����U  ���justforfun_justforfun_ ���U  �����U  P����U  �����U  @����U  �|g��+n��1&/      Some_stuffs �����U  �����U  ���justforfun_justforfun_ ���U  �����U  @����U  �����U  @����U  �/���y�n�3/      Meeting     0���U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �/���y�nv�3/       Workout     ���U  ���U  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   '��U  �/���y�nr�3/       Meeting     0 ��U  � ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �! ��U  a��H�C�p
"C/       Appointment  v��U  �v��U  `wjustforfun_justforfun_ ��U  �y��U  �z��U  `{��U  �{��U  b��H�C�p�!C/       Some_stuffs �M��U  �N��U  `OSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �T��U  c��H�C�p�(C/       Birthday    п��U  P���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  hR>Vs�qmc~&/      Birthday U  �� ��U  `� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0� ��U  ��-J/r��S/       Appointment �s��U  `t��U  �tSome_stuffs_Some_stuffs_ �U  `w��U  �w��U  �x��U  `y��U  ��-J/r�S/      Appointment ���U  p��U  0Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ���U  ��-J/r*�S/       Workout     p� ��U  0� ��U  �� justforfun_justforfun_  ��U  �� ��U  0� ��U  м ��U  �� ��U  �u�s#,uT<q/       Some_stuffs ���U  ����U  `�This_stuffs_This_stuffs_ �U   ���U  ���U  ����U   ���U  �u�s#,uT?q/       Appointment ����U   ���U  ��Some_stuffs_Some_stuffs_ �U  ����U  ����U  0���U  Щ��U  �u�s#,uO<q/       Appointment P���U  ����U  ��justforfun_justforfun_ ��U  P���U  ���U  ����U  ����U  �emvu�$t/       Workout ffs ����U  ���U  ЅThis_stuffs_This_stuffs_ �U  @���U  ����U  `���U  ����U  �emvu�$t/      Appointment ����U  0���U  �justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  ����U  �emvuE!t/       Meeting     `���U   ���U  ��Some_stuffs_Some_stuffs_ �U  ����U  p���U  ����U  ����U  ��-��vO�/      Workout ffs ����U  `���U  �justforfun_justforfun_ _This_stuffs_This_stuffs_ �U  ���U  ��-��v��/       Workout      &��U  �&��U  `'Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  p+��U  ��-��v��/       Appointment ����U  @���U  ��Some_stuffs_Some_stuffs_ �U  ���U  ����U  ���U  ����U  Y[����vEd�/       Appointment @� ��U   � ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   ��U  Z[����v�e�/       Some_stuffs ���U   '��U  PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �"��U  [[����v�h�/       Some_stuffs `_ ��U   ` ��U  `d This_stuffs_This_stuffs_ �U  �n ��U  Po ��U  �t ��U  �v ��U  ѣ��$*w���/      Birthday    г��U  ����U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  й��U  ң��$*w��/       Workout     �� ��U  `� ��U  �� This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �� ��U  ӣ��$*w��/       Birthday U  �U��U  pV��U  �Vjustforfun_justforfun_ ��U   Y��U  �Y��U  @Z��U   [��U  e��p�hx�G�/       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             e��p�hx�A�/       Meeting �U  � ��U  � ��U  � This_stuffs_This_stuffs_ �U   ! ��U  �! ��U  P% ��U  & ��U  e��p�hx�G�/       Some_stuffs �����U  �����U  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  @����U  ٶ�z��xT�/       Meeting �U  ����U  ���U  гSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  P���U  ڶ�z��xV�/       Some_stuffs  ��U  ���U  �This_stuffs_This_stuffs_ �U   ��U  ���U  `��U  ���U  ۶�z��xiZ�/       Appointment  ���U  ����U    This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  �G���@y7[ /       Appointment �� ��U  p� ��U  0� Some_stuffs_Some_stuffs_ �U   � ��U  �� ��U  �� ��U  @� ��U  �G���@y[ /       Some_stuffs �����U  �����U  ���This_stuffs_This_stuffs_ �U  �����U  @����U  �����U  @����U  �G���@y[ /       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_             �G���@y[ /      Birthday U  �M��U  �N��U  `OThis_stuffs_This_stuffs_ �U  �Q��U  �l��U  �S��U  �T��U  i����Uyi~&/       Workout �U   ���U  ����U  `�This_stuffs_This_stuffs_ �U  ���U  ����U  p���U  0���U  j����Uy]k~&/       Birthday    P����U  ����U  P��Some_stuffs_Some_stuffs_ �U  P����U  ����U  �����U  @����U  k����Uy e~&/       Appointment  ���U  ����U  `�This_stuffs_This_stuffs_ �U  ����U  @���U  ����U  p���U  l����Uyk~&/       Some_stuffs px��U  �x��U  pySome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  0}��U  m����Uy�k~&/       Meeting     ���U  ����U  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ���U  ��Cck�|���/      Some_stuffs �����U  `����U  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ��Cck�|g��/       Workout ffs  ���U  ����U   �justforfun_justforfun_ _This_stuffs_This_stuffs_ �U   ���U  ��Cck�|��/       Appointment P� ��U  � ��U  п This_stuffs_This_stuffs_ �U  �� ��U  �� ��U  P� ��U  �� ��U  �)o�_}z�/      Workout                        justforfun_justforfun_                                       �����6* /       Some_stuffs � ��U  � ��U  � This_stuffs_This_stuffs_ �U  0 ��U  � ��U  � ��U  � ��U  м��2��ڙ+ /       Some_stuffs � ��U  � ��U  � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  & ��U  �C���N�b&/       Meeting     ���U  ����U  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  �C���N��&/      Workout     м ��U  �� ��U  P� This_stuffs_This_stuffs_ �U  P� ��U  � ��U  �� ��U  �� ��U  �C���N�B&/       Workout     �`��U  Pa��U  �ajustforfun_justforfun_ _ �U  �c��U  Pd��U  �d��U  �e��U  ��Ga��&/      Birthday U  �7 ��U  �8 ��U  @< justforfun_justforfun_  ��U  pE ��U  0F ��U   J ��U  �J ��U  ��	���1&/       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_             aw��.�&/       Birthday    @� ��U   � ��U  �� This_stuffs_This_stuffs_ �U  � ��U  �� ��U  �� ��U  P� ��U  aw��!�&/       Some_stuffs  ��U  ���U  �This_stuffs_This_stuffs_ ome_stuffs_Some_stuffs_ �U  0��U  aw����&/       Birthday fs  p��U  �p��U   qThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  pu��U  aw����&/       Workout     �� ��U  �� ��U   � This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  `� ��U  = ��0*�j�[&/       Appointment �L��U  `M��U   NSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �R��U  = ��0*���[&/       Workout      <��U  �<��U  `>Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  `C��U  = ��0*���[&/      Some_stuffs `2��U   3��U  �3Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �8��U  Y��܆ת�jl&/       Some_stuffs ����U  `���U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   ��U  Z��܆ת�gl&/       Meeting     �l��U  Pm��U  �mjustforfun_justforfun_ _ �U  �~��U   ��U  �p��U  �q��U  [��܆ת%dl&/       Appointment �P��U  �Q��U  RSome_stuffs_Some_stuffs_ �U  PT��U  �T��U  PU��U  �U��U  ȁ�V����n&/       Meeting     p� ��U  0� ��U  �� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �� ��U  d�:�`b�!�{&/       Workout     p\��U  0]��U  �]This_stuffs_This_stuffs_ �U  �`��U  pa��U  0b��U  �b��U  �14�&�[�u�&/       Birthday    ����U  ����U  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  �14�&�[�I�&/       Meeting     ���U  p���U  �Some_stuffs_Some_stuffs_ �U  0���U  ���U  ����U  p���U  �14�&�[�x�&/       Workout     �P��U  `Q��U   RSome_stuffs_Some_stuffs_ �U  �T��U  Pc��U  �V��U  �W��U  ����W�~�dy�&/      Meeting     ���U  0��U  �This_stuffs_This_stuffs_ �U  `��U   ��U  ���U  `��U  ¼��W�~�~�&/       Birthday    ����U  @���U   �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ����U  ü��W�~��}�&/       Some_stuffs `K��U   L��U  �LSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   Q��U  ����Nܷe7* /       Birthday     0��U  �0��U   =Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �5��U  ����Nܷ�;* /       Meeting      $��U  �$��U   %justforfun_justforfun_ ��U  `'��U  �'��U  �(��U  P)��U  ����Nܷ�6* /       Workout     �O��U  pP��U  �PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  0U��U  ����Nܷ�6* /       Meeting                        Some_stuffs_Some_stuffs_                                     ����Nܷ=* /      Appointment 06��U  �6��U  07justforfun_justforfun_ ��U  p9��U  0:��U  �:��U  0;��U  Y��NZ`���-$/       Birthday     =��U  �=��U  `2This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U   7��U  Z��NZ`��#)$/       Some_stuffs e��U  �e��U  fThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �j��U  [��NZ`��p.$/       Workout     �B��U  pC��U  ` Some_stuffs_Some_stuffs_ �U   #��U  �#��U   $��U  �$��U  \��NZ`���.$/       Birthday     v��U  �v��U   wThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  �{��U  ɑ�$����n&/      Appointment P��U  ��U  �This_stuffs_This_stuffs_ �U  �!��U  �"��U  P#��U  $��U  ʑ�$�Փ�n&/       Appointment �� ��U  �� ��U  P� Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U   � ��U  ˑ�$��|�n&/       Workout     ���U  @��U  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  ���U  ̑�$�Ւ�n&/       Birthday    ����U  @���U   �justforfun_justforfun_ _ �U  ����U  @���U  ����U  @���U  �)�	h��և	�/       Birthday    ����U  ����U  @�justforfun_justforfun_ ��U  ����U   ���U  ����U  @���U  �)�	h��֌�/       Appointment �Y��U  �Z��U  0[Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �_��U  �)�	h��֞�/       Appointment �� ��U  @� ��U  � This_stuffs_This_stuffs_ �U  �� ��U  P� ��U   � ��U  �� ��U  �)�	h�����/       Meeting     �F��U  @G��U  �GSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  �K��U  Q���~N�����&/       Workout     P����U  ����U  P��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ �U  @����U  R���~N����&/      Some_stuffs P����U  ����U  P��This_stuffs_This_stuffs_ �U  P����U  ����U  �����U  @����U  S���~N�۪��&/       Meeting     Pg��U  h��U  �hjustforfun_justforfun_ ��U  �k��U  l��U  �l��U  Pm��U  T���~N����&/       Birthday    ����U   ���U  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  U���~N�ۭ��&/       Appointment  ��U  ���U  �Some_stuffs_Some_stuffs_ �U  ���U  ���U  p��U  0��U  aOݱۭ��۳ /       Birthday    � ��U  � ��U  � Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  � ��U  bOݱۭ�޳ /       Birthday U  �E��U  0F��U  �FThis_stuffs_This_stuffs_ �U  �H��U  PI��U  J��U  �J��U  cOݱۭ��߳ /       Birthday    ����U  ����U   �justforfun_justforfun_ ��U   ���U  ����U  @���U   ���U  dOݱۭ�2س /       Appointment ���U  `���U  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ �U  ����U  