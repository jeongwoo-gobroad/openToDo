ܦ
 /   ��
 /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �< /   �< /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             8{ /   H{ /      Meeting                        This_stuffs_                                                                                                                                                                                                                                                         | /   � /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �lw /   -mw /       Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ,q /   ]q /      Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         \�; /   w�; /      Meeting                        justforfun                                                                                                                                                                                                                                                           }f /   >}f /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �c: /   �c: /      Workout                        This_stuffs_                                                                                                                                                                                                                                                         �|� /   /}� /   	   Workout                        This_stuffs_                                                                                                                                                                                                                                                         P� /   h� /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �G- /   �G- /      Meeting                        This_stuffs_                                                                                                                                                                                                                                                         � /   9� /      Some_stuffs                    This_stuffs_                                                                                                                                                                                                                                                         ��H /   ��H /      Some_stuffs                    justforfun                                                                                                                                                                                                                                                           l+� /   �+� /      Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         �p� /   #q� /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �= /   �= /      Meeting                        This_stuffs_                                                                                                                                                                                                                                                          9 /   K9 /      Workout                        This_stuffs_                                                                                                                                                                                                                                                         4�V /   G�V /      Birthday                       This_stuffs_                                                                                                                                                                                                                                                         �Ǵ /   �Ǵ /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             4� /   g� /       Birthday                       justforfun                                                                                                                                                                                                                                                           D�v /   o�v /       Workout                        This_stuffs_                                                                                                                                                                                                                                                         �y /   (�y /      Workout                        justforfun                                                                                                                                                                                                                                                           X' /   p' /      Birthday                       justforfun                                                                                                                                                                                                                                                           ;< /   A;< /      Birthday                       justforfun                                                                                                                                                                                                                                                           � /   '� /      Appointment                    Some_stuffs_                                                                                                                                                                                                                                                         -q /   ^v /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �|� /   �z� /       Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         �z� /   �z� /       Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ؓ� /   ٓ� /       Some_stuffs                    This_stuffs_                                                                                                                                                                                                                                                         lqZ /   uqZ /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             t� /   u� /   	   Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��� /   ��� /      Birthday                       Some_stuffs_                                                                                                                                                                                                                                                         <�f /   \�f /      Workout                        justforfun                                                                                                                                                                                                                                                           �X /   �X /   	   Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             P� /   }� /       Some_stuffs                    justforfun                                                                                                                                                                                                                                                           N� /   $N� /      Appointment                    justforfun                                                                                                                                                                                                                                                           �[, /   �[, /      Birthday                       This_stuffs_                                                                                                                                                                                                                                                         ��J /   ��J /   	   Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��
 /   ��
 /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �r+ /   s+ /      Workout �U   %�N�U  p'�N�U  0)�This_stuffs_This_stuffs_ �U   2�N�U  �3�N�U  �6�N�U   8�N�U  ;�N�U  �<�N�U  �>�N�U   @�N�U  @B�N�U  �D�N�U  H�N�U  �I�N�U  �K�N�U  PM�N�U  �O�N�U   Q�N�U  �S�N�U  �T�N�U  �V�N�U  pX�N�U   \�N�U  �]�N�U  `�N�U  �b�N�U  @e�N�U  �f�N�U  pi�N�U  �j�N�U  �m�N�U  �;i /   �;i /      Workout                        Some_stuffs_                                                                                                                                                                                                                                                         ��� /   N�� /       Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �Г /   �Г /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             \D� /   fD� /      Meeting                        justforfun                                                                                                                                                                                                                                                            �+ /   "�+ /      Appointment                    This_stuffs_                                                                                                                                                                                                                                                         �Ǵ /   CŴ /      Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         @T� /   GT� /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �*� /   �*� /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             _I /   J_I /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �TK /   �TK /       Appointment                    This_stuffs_                                                                                                                                                                                                                                                         du; /   �u; /      Some_stuffs                    justforfun                                                                                                                                                                                                                                                           h� /   �� /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             `H+ /   wH+ /   	   Some_stuffs                    justforfun                                                                                                                                                                                                                                                           4� /   5� /   	   Some_stuffs                    This_stuffs_                                                                                                                                                                                                                                                         ��Z /   ��Z /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             8�w /   X�w /      Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         �(� /   �(� /       Some_stuffs                    justforfun                                                                                                                                                                                                                                                           xlg /   �lg /      Workout                        Some_stuffs_                                                                                                                                                                                                                                                         �|� /   Pz� /      Workout                        This_stuffs_                                                                                                                                                                                                                                                         �lw /   �ow /      Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         8؆ /   V؆ /      Appointment                    justforfun                                                                                                                                                                                                                                                           �1 /   2 /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             4�� /   5�� /      Meeting                        This_stuffs_                                                                                                                                                                                                                                                         !9 /   9 /      Birthday                       Some_stuffs_                                                                                                                                                                                                                                                         4� /   :� /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �x /   �x /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��� /   ��� /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �lw /   �nw /   	   Some_stuffs                    justforfun                                                                                                                                                                                                                                                           �X /   �X /      Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         H�� /   {�� /   	   Workout                        Some_stuffs_                                                                                                                                                                                                                                                         |?� /   ~?� /      Meeting                        justforfun                                                                                                                                                                                                                                                           `MX /   `MX /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             u� /   Iu� /      Meeting                        Some_stuffs_                                                                                                                                                                                                                                                         �: /   �: /      Birthday                       justforfun                                                                                                                                                                                                                                                           m+� /   �(� /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �Y /   �Y /      Workout                        This_stuffs_                                                                                                                                                                                                                                                         <~
 /   d~
 /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �� /   �� /      Workout                        justforfun                                                                                                                                                                                                                                                           5� /   $� /      Birthday                       justforfun                                                                                                                                                                                                                                                           <@W /   N@W /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �x /   Bx /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��� /   ��� /      Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         �, /   9�, /       Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �-� /   �-� /      Appointment                    This_stuffs_                                                                                                                                                                                                                                                         �1 /   . /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             � /   � /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �c: /   �f: /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��* /   ��* /      Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         d� /   Fd� /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             xO /   �O /      Workout                        This_stuffs_                                                                                                                                                                                                                                                         �r- /   �r- /      Appointment                    justforfun                                                                                                                                                                                                                                                           �m� /   �m� /      Some_stuffs                    Some_stuffs_                                                                                                                                                                                                                                                         \�+ /   ��+ /      Birthday                       This_stuffs_                                                                                                                                                                                                                                                         ��g /   ɳg /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �p� /   dx� /      Appointment                    justforfun                                                                                                                                                                                                                                                           �{h /   %|h /      Workout                        Some_stuffs_                                                                                                                                                                                                                                                         �G /   D�G /      Appointment                    Some_stuffs_                                                                                                                                                                                                                                                         �$+ /   %+ /   	   Meeting                        Some_stuffs_                                                                                                                                                                                                                                                         ��, /   ��, /       Meeting                        This_stuffs_                                                                                                                                                                                                                                                          �; /   $�; /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                              �K /   <�K /       Birthday                       justforfun                                                                                                                                                                                                                                                           �+ /   "�+ /   	   Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             d� /   �� /      Birthday                       justforfun                                                                                                                                                                                                                                                           0x� /   Kx� /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             u� /   6� /      Birthday                       justforfun                                                                                                                                                                                                                                                           � /   �� /   	   Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �˕ /   *̕ /      Meeting                        This_stuffs_                                                                                                                                                                                                                                                         ��� /   ʷ� /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��g /   ��g /      Appointment                    justforfun                                                                                                                                                                                                                                                           Ԕ� /   Ք� /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             D�Z /   _�Z /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             TPu /   �Pu /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �(� /   '� /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ࡗ /   �� /       Appointment                    Some_stuffs_                                                                                                                                                                                                                                                         �h /   �h /      Birthday                       Some_stuffs_                                                                                                                                                                                                                                                         �
f /   �
f /      Birthday                       Some_stuffs_                                                                                                                                                                                                                                                         P�K /   _�K /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ylg /   Hhg /       Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �$+ /   a#+ /      Meeting                        Some_stuffs_                                                                                                                                                                                                                                                         �m� /   �i� /      Workout                        justforfun                                                                                                                                                                                                                                                           �[ /   �[ /   	   Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �{h /   Mwh /      Meeting                        Some_stuffs_                                                                                                                                                                                                                                                         �?8 /   �?8 /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ̌W /   όW /       Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �� /   �� /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��f /   ��f /       Appointment                    Some_stuffs_                                                                                                                                                                                                                                                         8}x /   :}x /      Meeting                        This_stuffs_                                                                                                                                                                                                                                                         �� /   P�� /   	   Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��Y /   ��Y /      Appointment                    justforfun                                                                                                                                                                                                                                                           ��Y /   `�Y /      Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             @�w /   C�w /      Birthday                       justforfun                                                                                                                                                                                                                                                           ��� /   K� /      Some_stuffs  %�N�U  p'�N�U  0)�justforfun   �-�N�U  /�N�U   2�N�U  �3�N�U  �6�N�U   8�N�U  ;�N�U  �<�N�U  �>�N�U   @�N�U  @B�N�U  �D�N�U  H�N�U  �I�N�U  �K�N�U  PM�N�U  �O�N�U   Q�N�U  �S�N�U  �T�N�U  �V�N�U  pX�N�U   \�N�U  �]�N�U  `�N�U  �b�N�U  @e�N�U  �f�N�U  pi�N�U  �j�N�U  �m�N�U  ha� /   ha� /      Meeting �U  Py�N�U  �z�N�U  �}�This_stuffs_This_stuffs_ �U  ���N�U  @��N�U  p��N�U  ���N�U  0��N�U  ���N�U   ��N�U  ���N�U  ���N�U  `��N�U  ���N�U  П�N�U  P��N�U  Ф�N�U  `��N�U  ���N�U  @��N�U  ���N�U  p��N�U  ���N�U  0��N�U  ���N�U  ���N�U   ��N�U  ���N�U  `äN�U  ǤN�U  �ȤN�U  �̤N�U  � /   6� /      Workout �U  ��N�U  P��N�U  ���justforfun   ���N�U   �N�U  ��N�U  @�N�U  ��N�U  p�N�U  0�N�U  p�N�U  @�N�U  ��N�U  `�N�U  ��N�U  �$�N�U  &�N�U  �*�N�U  P,�N�U  `1�N�U  �2�N�U  �7�N�U  @9�N�U  p>�N�U  �?�N�U  0E�N�U  pF�N�U  �K�N�U  �L�N�U   R�N�U  `S�N�U  �X�N�U  PZ�N�U  �_�N�U  ]�+ /   v�+ /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �p� /   �r� /      Meeting �U   %�N�U  p'�N�U  0)�Some_stuffs_Some_stuffs_ �U   2�N�U  �3�N�U  �6�N�U   8�N�U  ;�N�U  �<�N�U  �>�N�U   @�N�U  @B�N�U  �D�N�U  H�N�U  �I�N�U  �K�N�U  PM�N�U  �O�N�U   Q�N�U  �S�N�U  �T�N�U  �V�N�U  pX�N�U   \�N�U  �]�N�U  `�N�U  �b�N�U  @e�N�U  �f�N�U  pi�N�U  �j�N�U  �m�N�U  1x� /   �|� /      Some_stuffs Py�N�U  �z�N�U  �}�justforfun    ��N�U  ���N�U  ���N�U  @��N�U  p��N�U  ���N�U  0��N�U  ���N�U   ��N�U  ���N�U  ���N�U  `��N�U  ���N�U  П�N�U  P��N�U  Ф�N�U  `��N�U  ���N�U  @��N�U  ���N�U  p��N�U  ���N�U  0��N�U  ���N�U  ���N�U   ��N�U  ���N�U  `äN�U  ǤN�U  �ȤN�U  �̤N�U  �&X /   �&X /      Birthday U  �ܤN�U  pޤN�U  p�Some_stuffs_  �N�U  ��N�U  ��N�U  `�N�U  ��N�U  P��N�U  ���N�U  P��N�U  ���N�U   �N�U  ��N�U  @�N�U  ��N�U  p�N�U  0�N�U  p�N�U  @�N�U  ��N�U  `�N�U  ��N�U  �$�N�U  &�N�U  �*�N�U  P,�N�U  `1�N�U  �2�N�U  �7�N�U  @9�N�U  p>�N�U  �?�N�U  0E�N�U  L /   n /      Meeting                        This_stuffs_                                                                                                                                                                                                                                                         � X /   � X /      Appointment  %�N�U  p'�N�U  0)�justforfun   �-�N�U  /�N�U   2�N�U  �3�N�U  �6�N�U   8�N�U  ;�N�U  �<�N�U  �>�N�U   @�N�U  @B�N�U  �D�N�U  H�N�U  �I�N�U  �K�N�U  PM�N�U  �O�N�U   Q�N�U  �S�N�U  �T�N�U  �V�N�U  pX�N�U   \�N�U  �]�N�U  `�N�U  �b�N�U  @e�N�U  �f�N�U  pi�N�U  �j�N�U  �m�N�U  ,�f /   >�f /      Workout �U  p��N�U  ���N�U  0��justforfun    ��N�U  ���N�U  ���N�U  `��N�U  ���N�U  П�N�U  P��N�U  Ф�N�U  `��N�U  ���N�U  @��N�U  ���N�U  p��N�U  ���N�U  0��N�U  ���N�U  ���N�U   ��N�U  ���N�U  `äN�U  ǤN�U  �ȤN�U  �̤N�U  ΤN�U  �ѤN�U  `ӤN�U  @פN�U  �ؤN�U  �ܤN�U  pޤN�U  p�N�U  ��� /   ��� /   	   Appointment ��N�U  p�N�U  0�Some_stuffs_Some_stuffs_ �U  `�N�U  ��N�U  �$�N�U  &�N�U  �*�N�U  P,�N�U  `1�N�U  �2�N�U  �7�N�U  @9�N�U  p>�N�U  �?�N�U  0E�N�U  pF�N�U  �K�N�U  �L�N�U   R�N�U  `S�N�U  �X�N�U  PZ�N�U  �_�N�U  Pa�N�U  �f�N�U  `h�N�U   n�N�U  @o�N�U  �i�N�U   k�N�U  �l�N�U  \�; /   ��; /      Workout                        Some_stuffs_                                                                                                                                                                                                                                                         !�K /   �K /       Some_stuffs  %�N�U  p'�N�U  0)�This_stuffs_This_stuffs_ �U   2�N�U  �3�N�U  �6�N�U   8�N�U  ;�N�U  �<�N�U  �>�N�U   @�N�U  @B�N�U  �D�N�U  H�N�U  �I�N�U  �K�N�U  PM�N�U  �O�N�U   Q�N�U  �S�N�U  �T�N�U  �V�N�U  pX�N�U   \�N�U  �]�N�U  `�N�U  �b�N�U  @e�N�U  �f�N�U  pi�N�U  �j�N�U  �m�N�U  �� /   � /   	   Appointment Py�N�U  �z�N�U  �}�This_stuffs_This_stuffs_ �U  ���N�U  @��N�U  p��N�U  ���N�U  0��N�U  ���N�U   ��N�U  ���N�U  ���N�U  `��N�U  ���N�U  П�N�U  P��N�U  Ф�N�U  `��N�U  ���N�U  @��N�U  ���N�U  p��N�U  ���N�U  0��N�U  ���N�U  ���N�U   ��N�U  ���N�U  `äN�U  ǤN�U  �ȤN�U  �̤N�U  p' /   �' /      Meeting �U  ��N�U  P��N�U  ���This_stuffs_ ���N�U   �N�U  ��N�U  @�N�U  ��N�U  p�N�U  0�N�U  p�N�U  @�N�U  ��N�U  `�N�U  ��N�U  �$�N�U  &�N�U  �*�N�U  P,�N�U  `1�N�U  �2�N�U  �7�N�U  @9�N�U  p>�N�U  �?�N�U  0E�N�U  pF�N�U  �K�N�U  �L�N�U   R�N�U  `S�N�U  �X�N�U  PZ�N�U  �_�N�U  D�) /   J�) /      Meeting                        justforfun                                                                                                                                                                                                                                                           �uj /   �uj /       Workout �U   %�N�U  p'�N�U  0)�justforfun   �-�N�U  /�N�U   2�N�U  �3�N�U  �6�N�U   8�N�U  ;�N�U  �<�N�U  �>�N�U   @�N�U  @B�N�U  �D�N�U  H�N�U  �I�N�U  �K�N�U  PM�N�U  �O�N�U   Q�N�U  �S�N�U  �T�N�U  �V�N�U  pX�N�U   \�N�U  �]�N�U  `�N�U  �b�N�U  @e�N�U  �f�N�U  pi�N�U  �j�N�U  �m�N�U  ��u /   ��u /      Some_stuffs p��N�U  ���N�U  0��This_stuffs_This_stuffs_ �U  ���N�U  `��N�U  ���N�U  П�N�U  P��N�U  Ф�N�U  `��N�U  ���N�U  @��N�U  ���N�U  p��N�U  ���N�U  0��N�U  ���N�U  ���N�U   ��N�U  ���N�U  `äN�U  ǤN�U  �ȤN�U  �̤N�U  ΤN�U  �ѤN�U  `ӤN�U  @פN�U  �ؤN�U  �ܤN�U  pޤN�U  p�N�U  D9� /   x9� /       Birthday U  ��N�U  p�N�U  0�Some_stuffs_Some_stuffs_ �U  `�N�U  ��N�U  �$�N�U  &�N�U  �*�N�U  P,�N�U  `1�N�U  �2�N�U  �7�N�U  @9�N�U  p>�N�U  �?�N�U  0E�N�U  pF�N�U  �K�N�U  �L�N�U   R�N�U  `S�N�U  �X�N�U  PZ�N�U  �_�N�U  Pa�N�U  �f�N�U  `h�N�U   n�N�U  @o�N�U  �i�N�U   k�N�U  �l�N�U  �5v /   �5v /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             n+� /   �"� /       Meeting �U   %�N�U  p'�N�U  0)�This_stuffs_ �-�N�U  /�N�U   2�N�U  �3�N�U  �6�N�U   8�N�U  ;�N�U  �<�N�U  �>�N�U   @�N�U  @B�N�U  �D�N�U  H�N�U  �I�N�U  �K�N�U  PM�N�U  �O�N�U   Q�N�U  �S�N�U  �T�N�U  �V�N�U  pX�N�U   \�N�U  �]�N�U  `�N�U  �b�N�U  @e�N�U  �f�N�U  pi�N�U  �j�N�U  �m�N�U  ��w /   ��w /      Appointment Py�N�U  �z�N�U  �}�This_stuffs_  ��N�U  ���N�U  ���N�U  @��N�U  p��N�U  ���N�U  0��N�U  ���N�U   ��N�U  ���N�U  ���N�U  `��N�U  ���N�U  П�N�U  P��N�U  Ф�N�U  `��N�U  ���N�U  @��N�U  ���N�U  p��N�U  ���N�U  0��N�U  ���N�U  ���N�U   ��N�U  ���N�U  `äN�U  ǤN�U  �ȤN�U  �̤N�U  � /   $� /      Some_stuffs ��N�U  P��N�U  ���This_stuffs_This_stuffs_ �U  ��N�U  @�N�U  ��N�U  p�N�U  0�N�U  p�N�U  @�N�U  ��N�U  `�N�U  ��N�U  �$�N�U  &�N�U  �*�N�U  P,�N�U  `1�N�U  �2�N�U  �7�N�U  @9�N�U  p>�N�U  �?�N�U  0E�N�U  pF�N�U  �K�N�U  �L�N�U   R�N�U  `S�N�U  �X�N�U  PZ�N�U  �_�N�U  � /   � /       Some_stuffs                    justforfun                                                                                                                                                                                                                                                           h�� /   ��� /      Workout �U   %�N�U  p'�N�U  0)�This_stuffs_ �-�N�U  /�N�U   2�N�U  �3�N�U  �6�N�U   8�N�U  ;�N�U  �<�N�U  �>�N�U   @�N�U  @B�N�U  �D�N�U  H�N�U  �I�N�U  �K�N�U  PM�N�U  �O�N�U   Q�N�U  �S�N�U  �T�N�U  �V�N�U  pX�N�U   \�N�U  �]�N�U  `�N�U  �b�N�U  @e�N�U  �f�N�U  pi�N�U  �j�N�U  �m�N�U  ��W /   ɯW /       Workout �U  p��N�U  ���N�U  0��Some_stuffs_Some_stuffs_ �U  ���N�U  `��N�U  ���N�U  П�N�U  P��N�U  Ф�N�U  `��N�U  ���N�U  @��N�U  ���N�U  p��N�U  ���N�U  0��N�U  ���N�U  ���N�U   ��N�U  ���N�U  `äN�U  ǤN�U  �ȤN�U  �̤N�U  ΤN�U  �ѤN�U  `ӤN�U  @פN�U  �ؤN�U  �ܤN�U  pޤN�U  p�N�U   iJ /   LiJ /      Birthday U  ��N�U  p�N�U  0�This_stuffs_This_stuffs_ �U  `�N�U  ��N�U  �$�N�U  &�N�U  �*�N�U  P,�N�U  `1�N�U  �2�N�U  �7�N�U  @9�N�U  p>�N�U  �?�N�U  0E�N�U  pF�N�U  �K�N�U  �L�N�U   R�N�U  `S�N�U  �X�N�U  PZ�N�U  �_�N�U  Pa�N�U  �f�N�U  `h�N�U   n�N�U  @o�N�U  �i�N�U   k�N�U  �l�N�U  �h /   ��h /      Meeting                        This_stuffs_                                                                                                                                                                                                                                                         �� /   � /      Meeting �U   %�N�U  p'�N�U  0)�Some_stuffs_ �-�N�U  /�N�U   2�N�U  �3�N�U  �6�N�U   8�N�U  ;�N�U  �<�N�U  �>�N�U   @�N�U  @B�N�U  �D�N�U  H�N�U  �I�N�U  �K�N�U  PM�N�U  �O�N�U   Q�N�U  �S�N�U  �T�N�U  �V�N�U  pX�N�U   \�N�U  �]�N�U  `�N�U  �b�N�U  @e�N�U  �f�N�U  pi�N�U  �j�N�U  �m�N�U  �� /   �� /       Workout �U  p��N�U  ���N�U  0��justforfun    ��N�U  ���N�U  ���N�U  `��N�U  ���N�U  П�N�U  P��N�U  Ф�N�U  `��N�U  ���N�U  @��N�U  ���N�U  p��N�U  ���N�U  0��N�U  ���N�U  ���N�U   ��N�U  ���N�U  `äN�U  ǤN�U  �ȤN�U  �̤N�U  ΤN�U  �ѤN�U  `ӤN�U  @פN�U  �ؤN�U  �ܤN�U  pޤN�U  p�N�U  �� /   �� /      Some_stuffs ��N�U  p�N�U  0�Some_stuffs_Some_stuffs_ �U  `�N�U  ��N�U  �$�N�U  &�N�U  �*�N�U  P,�N�U  `1�N�U  �2�N�U  �7�N�U  @9�N�U  p>�N�U  �?�N�U  0E�N�U  pF�N�U  �K�N�U  �L�N�U   R�N�U  `S�N�U  �X�N�U  PZ�N�U  �_�N�U  Pa�N�U  �f�N�U  `h�N�U   n�N�U  @o�N�U  �i�N�U   k�N�U  �l�N�U  �Hw /   �Hw /      Meeting                        Some_stuffs_                                                                                                                                                                                                                                                         �r- /   �r- /      Some_stuffs  %�N�U  p'�N�U  0)�Some_stuffs_ �-�N�U  /�N�U   2�N�U  �3�N�U  �6�N�U   8�N�U  ;�N�U  �<�N�U  �>�N�U   @�N�U  @B�N�U  �D�N�U  H�N�U  �I�N�U  �K�N�U  PM�N�U  �O�N�U   Q�N�U  �S�N�U  �T�N�U  �V�N�U  pX�N�U   \�N�U  �]�N�U  `�N�U  �b�N�U  @e�N�U  �f�N�U  pi�N�U  �j�N�U  �m�N�U  �� /   W� /      Workout �U  Py�N�U  �z�N�U  �}�Some_stuffs_  ��N�U  ���N�U  ���N�U  @��N�U  p��N�U  ���N�U  0��N�U  ���N�U   ��N�U  ���N�U  ���N�U  `��N�U  ���N�U  П�N�U  P��N�U  Ф�N�U  `��N�U  ���N�U  @��N�U  ���N�U  p��N�U  ���N�U  0��N�U  ���N�U  ���N�U   ��N�U  ���N�U  `äN�U  ǤN�U  �ȤN�U  �̤N�U  �~ /   �~ /      Appointment �ܤN�U  pޤN�U  p�Some_stuffs_  �N�U  ��N�U  ��N�U  `�N�U  ��N�U  P��N�U  ���N�U  P��N�U  ���N�U   �N�U  ��N�U  @�N�U  ��N�U  p�N�U  0�N�U  p�N�U  @�N�U  ��N�U  `�N�U  ��N�U  �$�N�U  &�N�U  �*�N�U  P,�N�U  `1�N�U  �2�N�U  �7�N�U  @9�N�U  p>�N�U  �?�N�U  0E�N�U  &Z /   >&Z /      Workout �U  �f�N�U  `h�N�U   n�This_stuffs_This_stuffs_ �U  �l�N�U   u�N�U  �p�N�U   r�N�U  @s�N�U  �z�N�U  `v�N�U  �w�N�U  `y�N�U  ���N�U   |�N�U  @}�N�U  �~�N�U  ���N�U   ��N�U  ���N�U   ��N�U  ���N�U   ��N�U  @��N�U  ���N�U   ��N�U   ��N�U  ���N�U   ��N�U  @��N�U  @��N�U  ���N�U  @      �X /   J�X /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �Z� /   �Z� /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             I�� /   ݵ� /       Appointment  %�N�U  p'�N�U  0)�This_stuffs_This_stuffs_ �U   2�N�U  �3�N�U  �6�N�U   8�N�U  ;�N�U  �<�N�U  �>�N�U   @�N�U  @B�N�U  �D�N�U  H�N�U  �I�N�U  �K�N�U  PM�N�U  �O�N�U   Q�N�U  �S�N�U  �T�N�U  �V�N�U  pX�N�U   \�N�U  �]�N�U  `�N�U  �b�N�U  @e�N�U  �f�N�U  pi�N�U  �j�N�U  �m�N�U  yO /   �S /       Appointment Py�N�U  �z�N�U  �}�Some_stuffs_  ��N�U  ���N�U  ���N�U  @��N�U  p��N�U  ���N�U  0��N�U  ���N�U   ��N�U  ���N�U  ���N�U  `��N�U  ���N�U  П�N�U  P��N�U  Ф�N�U  `��N�U  ���N�U  @��N�U  ���N�U  p��N�U  ���N�U  0��N�U  ���N�U  ���N�U   ��N�U  ���N�U  `äN�U  ǤN�U  �ȤN�U  �̤N�U  $>� /   8>� /      Some_stuffs �ܤN�U  pޤN�U  p�This_stuffs_  �N�U  ��N�U  ��N�U  `�N�U  ��N�U  P��N�U  ���N�U  P��N�U  ���N�U   �N�U  ��N�U  @�N�U  ��N�U  p�N�U  0�N�U  p�N�U  @�N�U  ��N�U  `�N�U  ��N�U  �$�N�U  &�N�U  �*�N�U  P,�N�U  `1�N�U  �2�N�U  �7�N�U  @9�N�U  p>�N�U  �?�N�U  0E�N�U  �0h /   1h /      Workout �U  �i�N�U   k�N�U  �l�This_stuffs_ �p�N�U   r�N�U  @s�N�U  �z�N�U  `v�N�U  �w�N�U  `y�N�U  ���N�U   |�N�U  @}�N�U  �~�N�U  ���N�U   ��N�U  ���N�U   ��N�U  ���N�U   ��N�U  @��N�U  ���N�U   ��N�U   ��N�U  ���N�U   ��N�U  @��N�U  @��N�U  ���N�U  @��N�U  ���N�U  ���N�U  ���N�U   ��N�U  _I /   YI /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �� /   �� /      Workout                        Some_stuffs_                                                                                                                                                                                                                                                         �� /   R� /      Meeting �U   %�N�U  p'�N�U  0)�Some_stuffs_ �-�N�U  /�N�U   2�N�U  �3�N�U  �6�N�U   8�N�U  ;�N�U  �<�N�U  �>�N�U   @�N�U  @B�N�U  �D�N�U  H�N�U  �I�N�U  �K�N�U  PM�N�U  �O�N�U   Q�N�U  �S�N�U  �T�N�U  �V�N�U  pX�N�U   \�N�U  �]�N�U  `�N�U  �b�N�U  @e�N�U  �f�N�U  pi�N�U  �j�N�U  �m�N�U  \�� /   ~�� /      Appointment Py�N�U  �z�N�U  �}�Some_stuffs_  ��N�U  ���N�U  ���N�U  @��N�U  p��N�U  ���N�U  0��N�U  ���N�U   ��N�U  ���N�U  ���N�U  `��N�U  ���N�U  П�N�U  P��N�U  Ф�N�U  `��N�U  ���N�U  @��N�U  ���N�U  p��N�U  ���N�U  0��N�U  ���N�U  ���N�U   ��N�U  ���N�U  `äN�U  ǤN�U  �ȤN�U  �̤N�U  Pٳ /   lٳ /      Some_stuffs ��N�U  P��N�U  ���This_stuffs_ ���N�U   �N�U  ��N�U  @�N�U  ��N�U  p�N�U  0�N�U  p�N�U  @�N�U  ��N�U  `�N�U  ��N�U  �$�N�U  &�N�U  �*�N�U  P,�N�U  `1�N�U  �2�N�U  �7�N�U  @9�N�U  p>�N�U  �?�N�U  0E�N�U  pF�N�U  �K�N�U  �L�N�U   R�N�U  `S�N�U  �X�N�U  PZ�N�U  �_�N�U  	&Z /   �'Z /      Appointment `v�N�U  �w�N�U  `y�This_stuffs_  |�N�U  @}�N�U  �~�N�U  ���N�U   ��N�U  ���N�U   ��N�U  ���N�U   ��N�U  @��N�U  ���N�U   ��N�U   ��N�U  ���N�U   ��N�U  @��N�U  @��N�U  ���N�U  @��N�U  ���N�U  ���N�U  ���N�U   ��N�U  `��N�U  0��N�U  p��N�U  ࠥN�U   ��N�U  `��N�U  थN�U  @      ��: /   ܏: /   	   Some_stuffs                    This_stuffs_                                                                                                                                                                                                                                                         E�v /   ��v /      Appointment                    Some_stuffs_                                                                                                                                                                                                                                                         o+� /   �(� /      Some_stuffs  %�N�U  p'�N�U  0)�Some_stuffs_Some_stuffs_ �U   2�N�U  �3�N�U  �6�N�U   8�N�U  ;�N�U  �<�N�U  �>�N�U   @�N�U  @B�N�U  �D�N�U  H�N�U  �I�N�U  �K�N�U  PM�N�U  �O�N�U   Q�N�U  �S�N�U  �T�N�U  �V�N�U  pX�N�U   \�N�U  �]�N�U  `�N�U  �b�N�U  @e�N�U  �f�N�U  pi�N�U  �j�N�U  �m�N�U  �ky /   �ky /       Meeting     ���N�U  @��N�U  p��Some_stuffs_Some_stuffs_ �U   ��N�U  ���N�U  ���N�U  `��N�U  ���N�U  П�N�U  P��N�U  Ф�N�U  `��N�U  ���N�U  @��N�U  ���N�U  p��N�U  ���N�U  0��N�U  ���N�U  ���N�U   ��N�U  ���N�U  `äN�U  ǤN�U  �ȤN�U  �̤N�U  ΤN�U  �ѤN�U  `ӤN�U  @פN�U  �ؤN�U  �ܤN�U  �� /   �� /      Meeting �U  ���N�U  P��N�U  ���Some_stuffs_ ��N�U  @�N�U  ��N�U  p�N�U  0�N�U  p�N�U  @�N�U  ��N�U  `�N�U  ��N�U  �$�N�U  &�N�U  �*�N�U  P,�N�U  `1�N�U  �2�N�U  �7�N�U  @9�N�U  p>�N�U  �?�N�U  0E�N�U  pF�N�U  �K�N�U  �L�N�U   R�N�U  `S�N�U  �X�N�U  PZ�N�U  �_�N�U  Pa�N�U  �f�N�U  AT� /   W� /       Workout �U  `y�N�U  ���N�U   |�justforfun   �~�N�U  ���N�U   ��N�U  ���N�U   ��N�U  ���N�U   ��N�U  @��N�U  ���N�U   ��N�U   ��N�U  ���N�U   ��N�U  @��N�U  @��N�U  ���N�U  @��N�U  ���N�U  ���N�U  ���N�U   ��N�U  `��N�U  0��N�U  p��N�U  ࠥN�U   ��N�U  `��N�U  थN�U  0��N�U  p��N�U  ���N�U  �� /   ¤ /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             i� /   � /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             <GZ /   cGZ /      Appointment  %�N�U  p'�N�U  0)�This_stuffs_ �-�N�U  /�N�U   2�N�U  �3�N�U  �6�N�U   8�N�U  ;�N�U  �<�N�U  �>�N�U   @�N�U  @B�N�U  �D�N�U  H�N�U  �I�N�U  �K�N�U  PM�N�U  �O�N�U   Q�N�U  �S�N�U  �T�N�U  �V�N�U  pX�N�U   \�N�U  �]�N�U  `�N�U  �b�N�U  @e�N�U  �f�N�U  pi�N�U  �j�N�U  �m�N�U  �[ /   �[ /      Some_stuffs p��N�U  ���N�U  0��justforfun    ��N�U  ���N�U  ���N�U  `��N�U  ���N�U  П�N�U  P��N�U  Ф�N�U  `��N�U  ���N�U  @��N�U  ���N�U  p��N�U  ���N�U  0��N�U  ���N�U  ���N�U   ��N�U  ���N�U  `äN�U  ǤN�U  �ȤN�U  �̤N�U  ΤN�U  �ѤN�U  `ӤN�U  @פN�U  �ؤN�U  �ܤN�U  pޤN�U  p�N�U  L�h /   �h /       Some_stuffs ��N�U  p�N�U  0�This_stuffs_ @�N�U  ��N�U  `�N�U  ��N�U  �$�N�U  &�N�U  �*�N�U  P,�N�U  `1�N�U  �2�N�U  �7�N�U  @9�N�U  p>�N�U  �?�N�U  0E�N�U  pF�N�U  �K�N�U  �L�N�U   R�N�U  `S�N�U  �X�N�U  PZ�N�U  �_�N�U  Pa�N�U  �f�N�U  `h�N�U   n�N�U  @o�N�U  �i�N�U   k�N�U  �l�N�U  @b� /   ub� /      Meeting �U   ��N�U  ���N�U   ��This_stuffs_This_stuffs_ �U  ���N�U   ��N�U   ��N�U  ���N�U   ��N�U  @��N�U  @��N�U  ���N�U  @��N�U  ���N�U  ���N�U  ���N�U   ��N�U  `��N�U  0��N�U  p��N�U  ࠥN�U   ��N�U  `��N�U  थN�U  0��N�U  p��N�U  ���N�U  �N�U  p��N�U  �N�U  ���N�U   ��N�U  �N�U  �^� /   �^� /      Meeting �U   %�N�U  p'�N�U  0)�This_stuffs_This_stuffs_ �U   2�N�U  �3�N�U  �6�N�U   8�N�U  ;�N�U  �<�N�U  �>�N�U   @�N�U  @B�N�U  �D�N�U  H�N�U  �I�N�U  �K�N�U  PM�N�U  �O�N�U   Q�N�U  �S�N�U  �T�N�U  �V�N�U  pX�N�U   \�N�U  �]�N�U  `�N�U  �b�N�U  @e�N�U  �f�N�U  pi�N�U  �j�N�U  �m�N�U   /   E /      Appointment p��N�U  ���N�U  0��This_stuffs_  ��N�U  ���N�U  ���N�U  `��N�U  ���N�U  П�N�U  P��N�U  Ф�N�U  `��N�U  ���N�U  @��N�U  ���N�U  p��N�U  ���N�U  0��N�U  ���N�U  ���N�U   ��N�U  ���N�U  `äN�U  ǤN�U  �ȤN�U  �̤N�U  ΤN�U  �ѤN�U  `ӤN�U  @פN�U  �ؤN�U  �ܤN�U  pޤN�U  p�N�U  �H /    �H /      Appointment ��N�U  p�N�U  0�This_stuffs_ @�N�U  ��N�U  `�N�U  ��N�U  �$�N�U  &�N�U  �*�N�U  P,�N�U  `1�N�U  �2�N�U  �7�N�U  @9�N�U  p>�N�U  �?�N�U  0E�N�U  pF�N�U  �K�N�U  �L�N�U   R�N�U  `S�N�U  �X�N�U  PZ�N�U  �_�N�U  Pa�N�U  �f�N�U  `h�N�U   n�N�U  @o�N�U  �i�N�U   k�N�U  �l�N�U  �G /   x�G /      Appointment  ��N�U  ���N�U   ��This_stuffs_This_stuffs_ �U  ���N�U   ��N�U   ��N�U  ���N�U   ��N�U  @��N�U  @��N�U  ���N�U  @��N�U  ���N�U  ���N�U  ���N�U   ��N�U  `��N�U  0��N�U  p��N�U  ࠥN�U   ��N�U  `��N�U  थN�U  0��N�U  p��N�U  ���N�U  �N�U  p��N�U  �N�U  ���N�U   ��N�U  �N�U  |�* /   ��* /      Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��8 /   ��8 /      Meeting                        justforfun                                                                                                                                                                                                                                                           � /   � /   	   Appointment  %�N�U  p'�N�U  0)�justforfun   �-�N�U  /�N�U   2�N�U  �3�N�U  �6�N�U   8�N�U  ;�N�U  �<�N�U  �>�N�U   @�N�U  @B�N�U  �D�N�U  H�N�U  �I�N�U  �K�N�U  PM�N�U  �O�N�U   Q�N�U  �S�N�U  �T�N�U  �V�N�U  pX�N�U   \�N�U  �]�N�U  `�N�U  �b�N�U  @e�N�U  �f�N�U  pi�N�U  �j�N�U  �m�N�U  ]�� /   4�� /      Some_stuffs Py�N�U  �z�N�U  �}�This_stuffs_This_stuffs_ �U  ���N�U  @��N�U  p��N�U  ���N�U  0��N�U  ���N�U   ��N�U  ���N�U  ���N�U  `��N�U  ���N�U  П�N�U  P��N�U  Ф�N�U  `��N�U  ���N�U  @��N�U  ���N�U  p��N�U  ���N�U  0��N�U  ���N�U  ���N�U   ��N�U  ���N�U  `äN�U  ǤN�U  �ȤN�U  �̤N�U  