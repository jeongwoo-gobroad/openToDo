>~
 /   �}
 /      Appointment �z�/V  ���/V  �~This_stuffs_This_stuffs_ /V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  ݦ
 /   ��
 /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ��
 /   k�
 /      Some_stuffs ���/V  ���/V  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V  $ /   [ /      Birthday     ��/V  @��/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  C /   6C /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �� /   $� /      Some_stuffs ��ӿ&V  P�ӿ&V  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  �� /   �� /      Birthday    �		�/V  �
	�/V  	Some_stuffs_Some_stuffs_ /V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  �� /   R� /      Meeting &V   �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  O /   n /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             2) /   k) /      Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �S /   �O /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             9{ /   H{ /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             6� /   � /      Appointment �	�/V  P�	�/V  ��	This_stuffs_This_stuffs_ /V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  Ю	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  �� /   �� /      Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  
 /   � /      Appointment �T
�/V  pV
�/V  �W
This_stuffs_This_stuffs_ /V  �]
�/V  0_
�/V  p`
�/V  �a
�/V  �z
�/V  �{
�/V  Pf
�/V  �g
�/V  i
�/V  Pj
�/V  �k
�/V  �l
�/V  n
�/V  Po
�/V  �p
�/V  Pr
�/V  �s
�/V  u
�/V  �v
�/V  �w
�/V  y
�/V  �
�/V  0}
�/V  p~
�/V  �
�/V  ��
�/V  0�
�/V  p�
�/V  ��
�/V  �= /   �= /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �� /   �� /   	   Appointment ���/V   ��/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �/V  P�/V  ��/V  �/V  -� /   � /      Meeting /V   ��/V  `��/V  мSome_stuffs_Some_stuffs_ /V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  �� /   �� /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     � /   5� /   	   Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             [' /   p' /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �Q /   4N /      Workout     p��/V  0��/V  ��Some_stuffs_Some_stuffs_ /V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  p /   ]q /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �� /   �� /       Workout &V  p[ӿ&V  �\ӿ&V  0`�justforfun_justforfun_ ӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  �� /   � /      Birthday V  �ӿ&V  p�ӿ&V  p��justforfun_justforfun_ ӿ&V  �ӿ&V  `�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  %� /   �� /      Workout /V  @	�/V  �,	�/V  �	justforfun_justforfun_ 	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  �[ /   �[ /   	   Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �~ /   �~ /      Appointment �ӿ&V  p�ӿ&V  p��Some_stuffs_Some_stuffs_ &V  �ӿ&V  `�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  � /   � /   	   Appointment ��/V  p�/V  pjustforfun_justforfun_ �/V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  � /   '� /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             5� /   :� /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ~ /   f /      Workout /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �o /   �o /      Meeting     �R�/V  �S�/V  UThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  �� /   �� /      Appointment  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  r� /   � /      Meeting /V  ��	�/V  0�	�/V  p�	justforfun_justforfun_ 	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  �
�/V  �
�/V  ��	�/V  �	�/V  P 
�/V  �
�/V  
�/V  P
�/V  �
�/V  
�/V  �
�/V  

�/V  �
�/V  
�/V  �$
�/V  �%
�/V   
�/V  `
�/V  �
�/V  
�/V  P
�/V  �
�/V  P
�/V  � /   � /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �. /   2 /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �W /   �W /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �� /   ¤ /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     � /   '� /      Meeting     `��/V  ���/V  0�This_stuffs_This_stuffs_ /V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  �� /   �� /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                      /   Y /      Workout     P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  |D /   �D /      Appointment ���/V  Ъ�/V  P�justforfun_justforfun_ �/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V  Q� /   h� /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                      /   E /      Appointment p[ӿ&V  �\ӿ&V  0`�This_stuffs_This_stuffs_ &V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  r' /   K( /      Appointment  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ��( /   ��( /      Meeting     `��/V  ��/V  `�justforfun_justforfun_ �/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  `��/V  0��/V  p��/V  ���/V   ��/V  `��/V  ���/V  0��/V  u') /   �%) /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �t) /   �t) /      Workout     ���/V  ���/V  �Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  Н) /   ��) /      Birthday V  PZ	�/V  �[	�/V  `L	This_stuffs_This_stuffs_ /V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  E�) /   J�) /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               �* /   �* /      Some_stuffs ���/V  ���/V   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  �5* /   �5* /      Some_stuffs ��ӿ&V  P�ӿ&V  ���Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  _�* /   ��* /      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ��* /   ��* /       Workout     @��/V  ���/V  ��justforfun_justforfun_ �/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V  ��* /   ��* /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��* /   �+ /   	   Meeting /V  ��	�/V  ��	�/V   �	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  I#+ /   %+ /   	   Meeting /V   <�/V  �F�/V  @?Some_stuffs_Some_stuffs_ /V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  aH+ /   wH+ /   	   Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               �r+ /   s+ /      Workout &V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �+ /   ڙ+ /       Some_stuffs � �/V  0�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  �+ /   "�+ /      Appointment  ��/V  @��/V  ��This_stuffs_This_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  G�+ /   ��+ /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ^, /   �[, /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �, /   �, /   	   Meeting     ���/V  ���/V   �justforfun_justforfun_ �/V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  ��, /   �, /      Birthday    ��/V  `�/V  �Some_stuffs_Some_stuffs_ /V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  �, /   9�, /       Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �G- /   �G- /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �r- /   Wq- /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �?8 /   �?8 /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �f8 /   0g8 /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��8 /   /�8 /      Appointment 0]�/V  p^�/V  �_justforfun_justforfun_ �/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  p9 /   K9 /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             h-9 /   p-9 /   	   Birthday    P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �W9 /   /R9 /      Appointment 0s�/V  pt�/V  �uSome_stuffs_Some_stuffs_ /V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  ��9 /   ��9 /      Meeting     ���/V   ��/V  @�justforfun_justforfun_ �/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  ��9 /   *�9 /      Workout     0]�/V  p^�/V  �_This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  �: /   �: /       Birthday     ��/V  @��/V  ��This_stuffs_This_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  �f: /   �c: /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��: /   ܏: /   	   Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                              �: /   '�: /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �(; /   /+; /      Meeting     ��/V  p�/V  pjustforfun_justforfun_ �/V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  \U; /   �U; /      Workout /V  �	�/V  P�	�/V  ��	This_stuffs_This_stuffs_ /V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  Ю	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  fu; /   �u; /      Appointment `��/V  ��/V  `�This_stuffs_This_stuffs_ /V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  `��/V  0��/V  p��/V  ���/V   ��/V  `��/V  ���/V  0��/V  ^�; /   ��; /      Appointment ���/V  Д�/V  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ��; /   $�; /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ]�; /   ��; /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �< /   �< /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ;< /   A;< /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �^< /   �f< /      Some_stuffs  <�/V  �F�/V  @?This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  -�< /   P�< /      Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             h�< /   ��< /      Appointment ��	�/V  Щ	�/V  �	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  XaG /   �aG /      Birthday V  `	�/V  �	�/V  	This_stuffs_This_stuffs_ /V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  ԨG /   �G /      Birthday    ���/V  0��/V  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  p�G /   D�G /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             iH /   �H /      Appointment ��ӿ&V  p�ӿ&V  0��This_stuffs_This_stuffs_ &V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  ��H /   ��H /      Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               <�H /    �H /      Appointment ��ӿ&V  p�ӿ&V  0��This_stuffs_This_stuffs_ &V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  �2I /   �2I /      Appointment ��/V  `�/V  �#This_stuffs_This_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  �XI /   J_I /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     p�I /   ��I /      Birthday    ���/V  ���/V   �This_stuffs_This_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  :�I /   ��I /       Some_stuffs ��/V  p�/V  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  ��I /   =�I /      Birthday    ��/V  P��/V  ��justforfun_justforfun_ �/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  �J /   -"J /      Meeting     �g	�/V  �h	�/V  P|	This_stuffs_This_stuffs_ /V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  "iJ /   poJ /      Appointment �
�/V  
�/V  P
justforfun_justforfun_ 
�/V  �
�/V  
�/V  P
�/V  � 
�/V  "
�/V  :
�/V   '
�/V  `(
�/V  �)
�/V  �*
�/V   ,
�/V  �-
�/V   /
�/V  `0
�/V  �1
�/V  `3
�/V  �4
�/V   6
�/V  �7
�/V  �N
�/V  P;
�/V  �<
�/V  >
�/V  �?
�/V  A
�/V  PB
�/V  �C
�/V  �D
�/V  F
�/V  ��J /   ��J /   	   Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     (�J /   <�J /      Appointment  ��/V  ���/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �TK /   �TK /       Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ؠK /   ڠK /      Birthday    �u	�/V  �v	�/V  `x	Some_stuffs_Some_stuffs_ /V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  |�K /   <�K /       Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               Q�K /   _�K /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     L�V /   l�V /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               p�V /   ��V /      Appointment @B�/V  �C�/V  PSome_stuffs_Some_stuffs_ /V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  6�V /   ��V /      Birthday    Ј�/V  P��/V  ЏThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  fW /   �W /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             >@W /   -AW /      Some_stuffs ���/V   ��/V  @�Some_stuffs_Some_stuffs_ /V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  paW /   �aW /      Workout     �!�/V  #�/V  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V  ͌W /   όW /       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ��W /   ɯW /       Workout &V  p[ӿ&V  �\ӿ&V  0`�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  P�W /   �W /      Meeting     �u	�/V  �v	�/V  `x	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��	�/V   �	�/V  @�	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  �X /   � X /      Appointment  �ҿ&V  p�ҿ&V  0��justforfun_justforfun_ ҿ&V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �&X /   �&X /      Birthday V  �ӿ&V  p�ӿ&V  p��Some_stuffs_Some_stuffs_ &V  �ӿ&V  `�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  aMX /   `MX /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     X�X /   �X /   	   Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ��X /   ��X /      Meeting     PZ	�/V  �[	�/V  `L	Some_stuffs_Some_stuffs_ /V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  ��X /   J�X /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �Y /   �Y /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �<Y /   �<Y /   	   Appointment ���/V   ��/V  `�Some_stuffs_Some_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  �Y /   ��Y /      Meeting     Ј�/V  P��/V  ЏSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  K�Y /   ��Y /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               �'Z /   >&Z /      Workout &V  �6Կ&V  `8Կ&V   >�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   BԿ&V  @CԿ&V  �JԿ&V  `FԿ&V  �GԿ&V  `IԿ&V  �PԿ&V   LԿ&V  @MԿ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @      ?GZ /   cGZ /      Appointment  �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  mqZ /   uqZ /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �Z /   _�Z /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ��Z /   ��Z /      Meeting     �R�/V  �S�/V  UThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  d	[ /   �[ /      Some_stuffs p[ӿ&V  �\ӿ&V  0`�justforfun_justforfun_ ӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  h	f /   �
f /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ?1f /   Q1f /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     }f /   {}f /      Workout /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ��f /   ��f /       Appointment ���/V   ��/V  `�Some_stuffs_Some_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  /�f /   >�f /      Workout &V  p[ӿ&V  �\ӿ&V  0`�justforfun_justforfun_ ӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  =�f /   \�f /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               Xg /   �g /   	   Some_stuffs �		�/V  �
	�/V  	This_stuffs_This_stuffs_ /V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  HBg /   {Bg /      Birthday V  T	�/V  PU	�/V  �V	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  /hg /   �lg /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             1�g /   ��g /      Some_stuffs P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��g /   ɳg /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ��g /   ��g /      Meeting     p[ӿ&V  �\ӿ&V  0`�This_stuffs_This_stuffs_ &V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  h /   h /      Meeting /V  `	�/V  �	�/V  	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  �0h /   1h /      Workout &V  �9Կ&V   ;Կ&V  �<�This_stuffs_This_stuffs_ &V  @CԿ&V  �JԿ&V  `FԿ&V  �GԿ&V  `IԿ&V  �PԿ&V   LԿ&V  @MԿ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  xh /   %|h /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��h /   �h /      Appointment @3	�/V  �4	�/V  �5	Some_stuffs_Some_stuffs_ /V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  [�h /   �h /       Some_stuffs ��ӿ&V  p�ӿ&V  0��This_stuffs_This_stuffs_ &V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  ��h /   �h /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �;i /   �;i /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             gi /   gi /      Appointment  ��/V  ���/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  ��i /   ��i /      Meeting     Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  t�i /   ~�i /      Appointment ���/V  Д�/V  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ��i /   �i /      Some_stuffs ���/V  Д�/V  �justforfun_justforfun_ �/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  QPj /   gPj /      Birthday V   �ҿ&V  p�ҿ&V  0��justforfun_justforfun_ ҿ&V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �uj /   �yj /      Appointment ��	�/V  0�	�/V  p�	Some_stuffs_Some_stuffs_ /V  ��	�/V  P�	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  0�	�/V  ��	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  �
�/V  �
�/V  ��	�/V  �	�/V  P 
�/V  �
�/V  
�/V  P
�/V  �
�/V  
�/V  �
�/V  

�/V  �
�/V  
�/V  �$
�/V  UPu /   �Pu /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ]pu /   Jou /      Some_stuffs �	�/V  P�	�/V  ��	Some_stuffs_Some_stuffs_ /V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  Ю	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��u /   ��u /      Some_stuffs p[ӿ&V  �\ӿ&V  0`�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  ��u /   ��u /       Some_stuffs ���/V  Д�/V  �justforfun_justforfun_ �/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ��u /   ��u /      Meeting     ��	�/V  Щ	�/V  �	justforfun_justforfun_ 	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  yv /   �v /   	   Appointment �Q	�/V  �R	�/V  T	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  �5v /   �8v /       Birthday    p��/V  ��/V  0�This_stuffs_This_stuffs_ /V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  p�/V  p�/V  _v /   1_v /      Appointment `	�/V  �	�/V  	Some_stuffs_Some_stuffs_ /V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  $�v /   K�v /      Workout /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  4�v /   X�v /      Appointment ���/V   ��/V  @�This_stuffs_This_stuffs_ /V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  �v /   o�v /       Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             w /   "w /      Birthday    � �/V  0�/V  pjustforfun_justforfun_ �/V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  �Hw /   �Hw /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �lw /   �nw /   	   Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               ��w /   0�w /   	   Appointment ���/V  0��/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  ��w /   C�w /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               :�w /   q�w /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             x /   �x /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     \^x /   �^x /      Birthday V  �	�/V  0�	�/V  p�	This_stuffs_This_stuffs_ /V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  p�	�/V  @�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V   �	�/V  `�	�/V  ��	�/V  P�	�/V  ��	�/V  0�	�/V  p�	�/V  9}x /   :}x /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �x /   �x /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��x /   �x /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               �y /   �y /      Some_stuffs ���/V   ��/V  `�justforfun_justforfun_ �/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  �ky /   �ky /       Meeting     �Vӿ&V  @Xӿ&V  p[�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  �y /   (�y /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               d� /   e� /      Appointment ���/V  ���/V   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  ��� /   ʷ� /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �� /   �� /      Some_stuffs �	�/V  P�	�/V  ��	justforfun_justforfun_ 	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  Ю	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V  �z� /   /}� /   	   Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             6�� /   ��� /       Meeting /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  � /   u� /   	   Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     }?� /   ~?� /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               Ab� /   ub� /      Meeting &V   RԿ&V  �SԿ&V   U�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  pԿ&V  �xԿ&V  �yԿ&V  p{Կ&V  �|Կ&V  ��Կ&V   �Կ&V  ��Կ&V  �� /   �� /      Birthday V   >Կ&V  @?Կ&V  �9�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �JԿ&V  `FԿ&V  �GԿ&V  `IԿ&V  �PԿ&V   LԿ&V  @MԿ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  9؆ /   V؆ /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               ��� /   ��� /   	   Appointment ��ӿ&V  p�ӿ&V  0��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  �"� /   �+� /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             IJ� /   �P� /      Appointment ��	�/V  ��	�/V   �	Some_stuffs_Some_stuffs_ /V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  �p� /   �r� /      Meeting &V   �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �� /   >�� /      Birthday    �	�/V  �/V  PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �� /   W� /       Birthday    PZ	�/V  �[	�/V  `L	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  � /   6� /      Workout &V  ��ӿ&V  P�ӿ&V  ���justforfun_justforfun_ ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  �;� /   �;� /      Appointment �#�/V  P%�/V  �)Some_stuffs_Some_stuffs_ /V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  �_� /   \_� /      Workout /V  �c
�/V  e
�/V  �O
This_stuffs_This_stuffs_ /V  �T
�/V  pV
�/V  �W
�/V  pY
�/V  �Z
�/V  0\
�/V  �]
�/V  0_
�/V  p`
�/V  �a
�/V  �z
�/V  �{
�/V  Pf
�/V  �g
�/V  i
�/V  Pj
�/V  �k
�/V  �l
�/V  n
�/V  Po
�/V  �p
�/V  Pr
�/V  �s
�/V  u
�/V  �v
�/V  �w
�/V  y
�/V  �
�/V  0}
�/V  g�� /   �� /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �؈ /   �؈ /   	   Meeting &V  �ӿ&V  p�ӿ&V  p��This_stuffs_This_stuffs_ &V  �ӿ&V  `�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  D�� /   ^�� /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     <Փ /   �Г /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     Q� /   }� /       Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               �E� /   �E� /      Some_stuffs T	�/V  PU	�/V  �V	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  �i� /   �m� /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ٓ� /   ٓ� /       Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             `� /   n� /      Workout     @��/V  � 	�/V  �	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  �-� /   n1� /      Meeting     P�/V  PQ�/V  0HSome_stuffs_Some_stuffs_ /V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  ��� /   ã� /   	   Birthday V  PZ	�/V  �[	�/V  `L	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �˕ /   
ʕ /      Appointment @��/V  � 	�/V  �	This_stuffs_This_stuffs_ /V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  �� /   �� /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �A� /   B� /      Workout     �#�/V  P%�/V  �)Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  �m� /   �m� /      Workout &V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  Ҳ� /   8�� /      Some_stuffs `��/V  ���/V  0�justforfun_justforfun_ �/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  �� /   � /      Birthday V  ��	�/V   �	�/V  @�	Some_stuffs_Some_stuffs_ /V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V   �	�/V  `�	�/V  ��	�/V  P�	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  0�	�/V  ��	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  �
�/V  �
�/V  ��	�/V  �	�/V  P 
�/V  Q� /   XR� /       Appointment ���/V   ��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  T~� /   W~� /       Appointment ��	�/V  ��	�/V   �	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  ڣ� /   �� /       Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             lŗ /   �ŗ /      Birthday    ���/V  P��/V  �This_stuffs_This_stuffs_ /V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V  �� /   �� /       Some_stuffs ���/V   ��/V  ��Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  �� /   �� /       Workout     P�/V  ��/V  This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  ;� /   p=� /      Birthday    ��ӿ&V  P�ӿ&V  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  �� /   �� /      Appointment ��/V  `�/V  �#This_stuffs_This_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  &>� /   �>� /      Meeting     ���/V  Ъ�/V  P�justforfun_justforfun_ �/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V  �a� /   �a� /      Some_stuffs ���/V  ���/V  �Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �� /   ~�� /      Appointment PIӿ&V  �Jӿ&V  �M�Some_stuffs_Some_stuffs_ &V  �Vӿ&V  @Xӿ&V  p[ӿ&V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  � /   �� /      Birthday V  �9Կ&V   ;Կ&V  �<�justforfun_justforfun_ Կ&V  @CԿ&V  �JԿ&V  `FԿ&V  �GԿ&V  `IԿ&V  �PԿ&V   LԿ&V  @MԿ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  Eף /   wף /      Workout &V   RԿ&V  �SԿ&V   U�Some_stuffs_Some_stuffs_ &V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  pԿ&V  �xԿ&V  �yԿ&V  p{Կ&V  �|Կ&V  ��Կ&V   �Կ&V  ��Կ&V  ��� /   4�� /      Some_stuffs  U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  %� /   �(� /       Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               1O� /   :O� /      Appointment p[ӿ&V  �\ӿ&V  0`�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  <o� /   Iu� /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             j�� /   ��� /       Some_stuffs Ј�/V  P��/V  ЏSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  E�� /   ��� /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �� /   �� /      Birthday V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V   8� /   "8� /      Birthday V  "
�/V  :
�/V   '
This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  `0
�/V  �1
�/V  `3
�/V  �4
�/V   6
�/V  �7
�/V  �N
�/V  P;
�/V  �<
�/V  >
�/V  �?
�/V  A
�/V  PB
�/V  �C
�/V  �D
�/V  F
�/V  PG
�/V  �H
�/V  �I
�/V  K
�/V  �L
�/V  �c
�/V  e
�/V  �O
�/V  0Q
�/V  pR
�/V  ia� /   ha� /      Meeting &V  PIӿ&V  �Jӿ&V  �M�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  Z�� /   �� /      Workout /V  �C
�/V  �D
�/V  F
Some_stuffs_Some_stuffs_ /V  K
�/V  �L
�/V  �c
�/V  e
�/V  �O
�/V  0Q
�/V  pR
�/V  �S
�/V  �T
�/V  pV
�/V  �W
�/V  pY
�/V  �Z
�/V  0\
�/V  �]
�/V  0_
�/V  p`
�/V  �a
�/V  �z
�/V  �{
�/V  Pf
�/V  �g
�/V  i
�/V  Pj
�/V  �k
�/V  �l
�/V  n
�/V  Po
�/V  �p
�/V  ��� /   ��� /      Birthday    P�/V  ��/V  Some_stuffs_Some_stuffs_ /V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  ]D� /   fD� /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               �k� /   �j� /       Appointment �z�/V  ���/V  �~Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ք� /   Ք� /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     %� /   �� /      Birthday    ���/V  @��/V  p�justforfun_justforfun_ �/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  �Z� /   �Z� /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �*� /   �*� /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     W� /   GT� /      Birthday V  ��/V  `�/V  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  �|� /   Kx� /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �� /   P�� /   	   Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �̲ /   Ͳ /      Workout &V  `sԿ&V  �tԿ&V  0~�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   �Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  @�Կ&V  @�Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  `�Կ&V  0�Կ&V  p�Կ&V   �Կ&V  @�Կ&V  ��Կ&V   �Կ&V  P�Կ&V  ��Կ&V  �Կ&V  0�Կ&V  p�Կ&V  ]�� /   � /      Meeting     � �/V  0�/V  pThis_stuffs_This_stuffs_ /V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  0@� /   X@� /       Birthday    �~�/V   ��/V  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  퍳 /   ��� /      Appointment ���/V  Д�/V  �justforfun_justforfun_ �/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ǵ� /   {�� /   	   Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ڳ /   lٳ /      Some_stuffs ��ӿ&V  P�ӿ&V  ���This_stuffs_This_stuffs_ &V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  �� /   �� /      Meeting &V  ��ӿ&V  P�ӿ&V  ���Some_stuffs_Some_stuffs_ &V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  N� /   $N� /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               �z� /   �z� /       Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �� /   7�� /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               CŴ /   �Ǵ /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     P� /   z� /      Workout     p�	�/V  ��	�/V  ��	justforfun_justforfun_ 	�/V   �	�/V  `�	�/V  ��	�/V  P�	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  0�	�/V  ��	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  �
�/V  �
�/V  ��	�/V  �	�/V  P 
�/V  �
�/V  
�/V  P
�/V  �
�/V  
�/V  �
�/V  

�/V  �
�/V  E9� /   x9� /       Birthday V  ��ӿ&V  p�ӿ&V  0��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  �^� /   �^� /      Meeting &V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  X�� /   n�� /      Some_stuffs �	�/V  0�	�/V  p�	Some_stuffs_Some_stuffs_ /V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  p�	�/V  @�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V   �	�/V  `�	�/V  ��	�/V  P�	�/V  ��	�/V  0�	�/V  p�	�/V  J�� /   1�� /      Some_stuffs ��/V  p�/V  pThis_stuffs_This_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  �Ե /   �Ե /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     (�� /   ��� /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     n$� /   �)� /      Appointment 0s�/V  pt�/V  �uThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  Hu� /   ou� /      Appointment `	�/V  �	�/V  	Some_stuffs_Some_stuffs_ /V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  ��� /   ��� /   	   Workout     ��/V  P��/V  ��This_stuffs_This_stuffs_ /V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ��� /   ��� /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             hrŭ}�  ��
 /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                      ���}�  H{ /      Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �+�}�  �= /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             x�j�}�  �� /      Meeting     ���/V  ���/V  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  ��p�}�  �� /       Workout                        justforfun_justforfun_                                                                                                                                                                                                                                                Ɲ�}�  V� /      Meeting /V  �
�/V  

�/V  �
justforfun_justforfun_ 
�/V   
�/V  `
�/V  �
�/V  
�/V  P
�/V  �
�/V  P
�/V  �
�/V  �
�/V  
�/V  P
�/V  � 
�/V  "
�/V  :
�/V   '
�/V  `(
�/V  �)
�/V  �*
�/V   ,
�/V  �-
�/V   /
�/V  `0
�/V  �1
�/V  `3
�/V  �4
�/V   6
�/V  �7
�/V  �N
�/V  P;
�/V   �A�}�  �[ /   	   Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     X��}�  �~ /      Appointment ���/V   ��/V  `�Some_stuffs_Some_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  ����}�  :� /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     P_i�}�  � /      Birthday    ���/V   ��/V  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  ���}�  ¤ /      Some_stuffs ��/V  `�/V  �#Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  �	�}�  A /      Appointment p��/V  ��/V  0�justforfun_justforfun_ �/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  p�/V  p�/V  ����}�  h� /      Birthday V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  x�� ~�  E /      Appointment @��/V  ���/V  ��This_stuffs_This_stuffs_ /V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  `��0~�  �') /       Birthday    �#�/V  P%�/V  �)This_stuffs_This_stuffs_ /V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  ��{3~�  J�) /      Meeting     �	�/V  �/V  Pjustforfun_justforfun_ �/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  В_5~�  �5* /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �9Z7~�  Ы* /      Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �~�7~�  ��* /      Some_stuffs `M�/V  �N�/V  �ZSome_stuffs_Some_stuffs_ /V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  XV�9~�  wH+ /   	   Some_stuffs Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  ���:~�  s+ /      Workout /V   <�/V  �F�/V  @?This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  8�:A~�  9�, /       Meeting     P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �-�q~�  �?8 /      Some_stuffs ���/V  @��/V  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  ��dv~�  �W9 /      Meeting     `	�/V  �	�/V  	This_stuffs_This_stuffs_ /V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  85�w~�  ��9 /       Some_stuffs ���/V   ��/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  ��{~�  ܏: /   	   Some_stuffs �W�/V  �X�/V  �eThis_stuffs_This_stuffs_ /V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  �n3~~�  �(; /      Appointment p`
�/V  �a
�/V  �z
justforfun_justforfun_ 
�/V  i
�/V  Pj
�/V  �k
�/V  �l
�/V  n
�/V  Po
�/V  �p
�/V  Pr
�/V  �s
�/V  u
�/V  �v
�/V  �w
�/V  y
�/V  �
�/V  0}
�/V  p~
�/V  �
�/V  ��
�/V  0�
�/V  p�
�/V  ��
�/V  ��
�/V  0�
�/V  ��
�/V  ��
�/V   �
�/V  ��
�/V   �
�/V  `�
�/V  �-x�~�  ��; /      Workout     P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��΂~�  A;< /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               ���~�  P�< /      Appointment ���/V  Д�/V  �This_stuffs_This_stuffs_ /V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ���~�  �H /      Appointment ���/V   ��/V  `�This_stuffs_This_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  @�̽~�  ��I /      Appointment ��	�/V  ��	�/V   �	Some_stuffs_Some_stuffs_ /V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  �|�~�  �J /       Appointment @	�/V  �,	�/V  �	Some_stuffs_Some_stuffs_ /V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  ��\�~�  ��J /   	   Meeting /V  ���/V  ���/V   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  XQ�~�  _�K /      Some_stuffs � �/V  0�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  H1�~�  όW /       Meeting     ��/V  `�/V  �#Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  0(��~�  �&X /      Birthday V  U�/V  PV�/V  �WSome_stuffs_Some_stuffs_ /V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  �xl�~�  `MX /      Meeting /V  �Z�/V  �[�/V  �RSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V  � �  (�Y /      Birthday    P�/V  ��/V  This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  8��  uqZ /      Meeting /V  ���/V   ��/V  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  �jw:�  \�f /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               �=�  2�g /      Some_stuffs P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  (�?>�  ��g /      Meeting      ��/V  @��/V  ��This_stuffs_This_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  pղ?�  1h /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �-D�  �;i /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �q�H�  gPj /      Birthday    ��/V  `�/V  �#justforfun_justforfun_ �/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  ��x�  �Pu /      Appointment  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �g�x�  �pu /      Meeting     p��/V  ��/V  0�Some_stuffs_Some_stuffs_ /V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  p�/V  p�/V  (�Ky�  ��u /      Some_stuffs �z�/V  ���/V  �~This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  �.X{�  �v /      Workout      ��/V  ���/V  ��This_stuffs_This_stuffs_ /V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  p���  :}x /      Meeting     �	�/V  �/V  PThis_stuffs_This_stuffs_ /V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �̺��  �ky /       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �S��  (�y /      Workout /V  ���/V  ���/V   �justforfun_justforfun_ �/V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  ЭE��  ʷ� /      Meeting /V  �W�/V  �X�/V  �eSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  �܄��  � /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               �����  ~?� /      Meeting /V  ��/V   �/V  �!justforfun_justforfun_ �/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  �n��  ub� /      Meeting     ���/V  0��/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  �}*��  �� /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     Ѕi��  V؆ /      Appointment Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  ���  ��� /   	   Appointment  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  8�S��  _J� /      Birthday    PZ	�/V  �[	�/V  `L	Some_stuffs_Some_stuffs_ /V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  ����  6� /      Workout     ��/V  `�/V  �#justforfun_justforfun_ �/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  H��  �؈ /   	   Meeting     ���/V   ��/V  `�This_stuffs_This_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  �Wj��  }� /       Some_stuffs P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  Hk��  ٓ� /       Some_stuffs  ��/V  @��/V  ��This_stuffs_This_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  �����  �� /      Meeting      ��/V  @��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ��_��  �m� /      Workout     ��/V  `�/V  �#This_stuffs_This_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P�e?��  �� /      Birthday    �	�/V  �/V  Pjustforfun_justforfun_ �/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  h�@��  wף /      Workout     �	�/V  �/V  PSome_stuffs_Some_stuffs_ /V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  ���@��  �� /      Some_stuffs "
�/V  :
�/V   '
Some_stuffs_Some_stuffs_ /V   ,
�/V  �-
�/V   /
�/V  `0
�/V  �1
�/V  `3
�/V  �4
�/V   6
�/V  �7
�/V  �N
�/V  P;
�/V  �<
�/V  >
�/V  �?
�/V  A
�/V  PB
�/V  �C
�/V  �D
�/V  F
�/V  PG
�/V  �H
�/V  �I
�/V  K
�/V  �L
�/V  �c
�/V  e
�/V  �O
�/V  0Q
�/V  pR
�/V  PiB��  :O� /      Appointment  ��/V  @��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���F��  ha� /      Meeting     ���/V  @��/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  `�mJ��  fD� /      Meeting     ��/V  `�/V  �#justforfun_justforfun_ �/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  �K��  l� /      Workout     P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ؂�K��  Ք� /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �O��  �Z� /      Appointment �z�/V  ���/V  �~Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  P��}��  �*� /      Birthday V  `M�/V  �N�/V  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  @      p?���  P�� /   	   Appointment P�/V  PQ�/V  0HThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  �H���  Ͳ /      Workout     0]�/V  p^�/V  �_This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  �N����  ��� /      Some_stuffs ���/V   ��/V  @�This_stuffs_This_stuffs_ /V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  `��/V  0��/V  p��/V  ���/V  訆���  #�� /      Workout     `M�/V  �N�/V  �ZSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  0|���  �� /      Meeting /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ������  $N� /      Appointment ��/V  p�/V  pjustforfun_justforfun_ �/V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  p����  �z� /       Workout     ��/V  `�/V  �#Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P۲���  x9� /       Birthday V  ���/V  P��/V  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V  ��S���  �^� /      Meeting /V   ��/V  `��/V  мThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  PVN���  �Ե /      Birthday    ��	�/V   �	�/V  p�	This_stuffs_This_stuffs_ /V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  p�	�/V  @�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ,?���  ��� /      Some_stuffs  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ���,�O d~
 /      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �R�-�O ��
 /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     x+�/�O _) /      Meeting &V  �(Կ&V  P*Կ&V  �/�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   ;Կ&V  �<Կ&V   EԿ&V  �@Կ&V   BԿ&V  @CԿ&V  �JԿ&V  `FԿ&V  �GԿ&V  `IԿ&V  �PԿ&V   LԿ&V  @MԿ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  ��]0�O g� /       Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               pL?/1�O  /      Workout     ���/V  ���/V   �This_stuffs_This_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  06EA3�O R /      Workout     �!�/V  #�/V  �Some_stuffs_Some_stuffs_ /V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V  P��H�O � /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �#�I�O �� /      Appointment ���/V   ��/V  ��Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  (��N�O �' /      Meeting &V  ��ӿ&V  P�ӿ&V  ���This_stuffs_This_stuffs_ &V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  ����d�O )�+ /   	   Birthday    ��/V   �/V  �!justforfun_justforfun_ �/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  h�ѭf�O ��, /       Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��{�O ��8 /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               H�.&}�O ��9 /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ���_}�O �: /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �|��O �u; /      Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               �n���O w�; /      Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               ���?��O �^< /      Birthday V   �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  P�S��O :�I /      Appointment ��Կ&V   �Կ&V  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  ��Կ&V  `�Կ&V  ��Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  `�Կ&V  0�Կ&V  p�Կ&V   �Կ&V  @�Կ&V  ��Կ&V   �Կ&V  P�Կ&V  ��Կ&V  �Կ&V  0�Կ&V  p�Կ&V  �Կ&V  `�Կ&V  ��Կ&V  ЩԿ&V  �Կ&V  P�Կ&V  ��Կ&V  �Կ&V  `ZA��O LiJ /      Birthday V  ��ӿ&V  p�ӿ&V  0��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  ���<��O G�V /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             (�6���O �W /      Meeting      <�/V  �F�/V  @?Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  0]�Ǯ�O N@W /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                      j���O ��Z /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     0a����O >}f /      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �V�P��O �uj /       Workout &V   �ҿ&V  p�ҿ&V  0��justforfun_justforfun_ ҿ&V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  nv���O �u /      Some_stuffs P�/V  ��/V  This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  h(7��O �5v /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �Z����O ��w /      Appointment PIӿ&V  �Jӿ&V  �M�This_stuffs_This_stuffs_ &V  �Vӿ&V  @Xӿ&V  p[ӿ&V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  @Rx��O X�w /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ��.<��O Fd� /      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     h=�L��O 5�� /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �FA3�O �� /   	   Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ����O �_� /       Appointment p[ӿ&V  �\ӿ&V  0`�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  ��*��O �-� /      Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �<��O *̕ /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �C	>�O 㲖 /      Meeting &V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  h����O � /   	   Appointment PIӿ&V  �Jӿ&V  �M�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  h�I�O Q� /      Birthday    ���/V  Ъ�/V  P�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V  �8C��O �� /      Workout &V  `FԿ&V  �GԿ&V  `I�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V   �&}/�O 8>� /      Some_stuffs �ӿ&V  p�ӿ&V  p��This_stuffs_This_stuffs_ &V  �ӿ&V  `�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  @�}�1�O ��� /      Workout &V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  ���X3�O f�� /      Appointment ��ӿ&V  p�ӿ&V  0��This_stuffs_This_stuffs_ &V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  �(��L�O �� /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               XJ��N�O K�� /      Birthday V  `FԿ&V  �GԿ&V  `I�Some_stuffs_Some_stuffs_ &V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  ��O�O �$� /      Meeting &V  `�Կ&V  ��Կ&V  `��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  p�Կ&V   �Կ&V  @�Կ&V  ��Կ&V   �Կ&V  P�Կ&V  ��Կ&V  �Կ&V  0�Կ&V  p�Կ&V  �Կ&V  `�Կ&V  ��Կ&V  ЩԿ&V  �Կ&V  P�Կ&V  ��Կ&V  �Կ&V  ��Կ&V  �Կ&V  `�Կ&V  ��Կ&V   �Կ&V  ��Կ&V  �Կ&V  �Կ&V  )1����� /       Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               *1����$� /      Some_stuffs ��/V  p�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  +1����� /       Some_stuffs Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  H�w2l��� /      Some_stuffs  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  x���3/� /   	   Some_stuffs  ��/V  @��/V  ��Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  �����F^v /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �����F]q /      Some_stuffs  ��/V  @��/V  ��Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  �����F^v /      Birthday V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �!��7� /      Birthday V  �9Կ&V   ;Կ&V  �<�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �GԿ&V  `IԿ&V  �PԿ&V   LԿ&V  @MԿ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  �!��7@� /      Birthday V   RԿ&V  �SԿ&V   U�justforfun_justforfun_ Կ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  pԿ&V  �xԿ&V  �yԿ&V  p{Կ&V  �|Կ&V  ��Կ&V   �Կ&V  ��Կ&V  �!��7� /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �!��7� /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �!��7@� /      Birthday    �	�/V  �/V  Pjustforfun_justforfun_ �/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �p�D�. /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �p�D�2 /      Appointment ���/V  ���/V   �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  �p�D�. /      Workout     Ј�/V  P��/V  ЏSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  ��t]�,	a#+ /      Meeting /V  �z�/V  ���/V  �~Some_stuffs_Some_stuffs_ /V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  ?��z�<	"�+ /   	   Meeting /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V   �Bh	�r- /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               a�&x��
9 /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             b�&x��
K9 /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             c�&x��
9 /      Birthday V   <�/V  �F�/V  @?Some_stuffs_Some_stuffs_ /V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  ��h}��
q�; /      Some_stuffs `FԿ&V  �GԿ&V  `I�justforfun_justforfun_ Կ&V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  ��h}��
$�; /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ��h}��
q�; /      Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               ��iHM,x�G /      Appointment  RԿ&V  �SԿ&V   U�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  pԿ&V  �xԿ&V  �yԿ&V  p{Կ&V  �|Կ&V  ��Կ&V   �Կ&V  ��Կ&V  ��iHM,D�G /      Appointment � �/V  0�/V  pSome_stuffs_Some_stuffs_ /V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  ��iHM,x�G /      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �5��0�)��H /   	   Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �5��0�) �H /      Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �5��0�)��H /   	   Meeting     P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  1����gx�K /       Some_stuffs  �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  2����gx<�K /       Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               3����gx�K /       Some_stuffs ��/V  p�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  i����X���W /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     j����X�� X /      Appointment ���/V  ���/V  �justforfun_justforfun_ �/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  k����X���W /      Meeting     p��/V  ���/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  �v�����X /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �v�����X /   	   Some_stuffs  U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �v�����X /      Some_stuffs ���/V   ��/V  ��Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  �x����J�X /      Workout     P�/V  PQ�/V  0HSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  �x������X /      Appointment  <�/V  �F�/V  @?Some_stuffs_Some_stuffs_ /V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  �x����5�X /      Appointment P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  q��0��[ /      Some_stuffs ��/V  `�/V  �justforfun_justforfun_ �/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  r��0�7[ /      Appointment P�/V  PQ�/V  0HSome_stuffs_Some_stuffs_ /V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  s��0�~[ /   	   Meeting     0��/V  ���/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V  �i�����f /   	   Meeting     �ӿ&V  p�ӿ&V  p��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  P�ӿ&V  ��ӿ&V  P�ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  �i�����
f /      Birthday    ���/V  ���/V   �Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  �i�����f /   	   Meeting     ���/V  `��/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  @�#U�s.ȣf /      Appointment @��/V  � 	�/V  �	justforfun_justforfun_ 	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  1�+�]Mwh /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             2�+�]%|h /      Workout     ���/V  ���/V   �Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  3�+�]Mwh /      Meeting /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ��l0�3j��h /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��l0�3j�h /      Birthday    Ј�/V  P��/V  ЏSome_stuffs_Some_stuffs_ /V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  ��l0�3j��h /      Meeting /V  �z�/V  ���/V  �~This_stuffs_This_stuffs_ /V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  h�K�T�-mw /       Some_stuffs ��/V  p�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  @��>����w /      Appointment P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ����E~#q� /      Birthday V  � �/V  0�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  ��S����ԓ /   	   Appointment  �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  ��S����Г /      Workout     ���/V  @��/V  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  ��S����ԓ /   	   Appointment ��/V  `�/V  �#This_stuffs_This_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  ��c��T4�� /      Some_stuffs PIӿ&V  �Jӿ&V  �M�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  ��c��T~�� /      Appointment @��/V  ���/V  `�Some_stuffs_Some_stuffs_ /V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  `��/V  0��/V  p��/V  ���/V   ��/V  `��/V  ��c��T4�� /      Some_stuffs Ј�/V  P��/V  ЏThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  ��&d'� /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ��&d�(� /       Some_stuffs                    justforfun_justforfun_                                                                                                                                                                                                                                               ��&d'� /      Birthday    P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ���kQo� /      Workout &V   �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  ���kIu� /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ���kQo� /      Workout /V  ���/V  P��/V  �Some_stuffs_Some_stuffs_ /V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V  pTp1,�sN�� /       Some_stuffs  U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ���۟w�� /      Birthday V  ��/V  P��/V  ��This_stuffs_This_stuffs_ /V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���۟w7� /      Workout     ��/V  p�/V  pThis_stuffs_This_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  ���۟w�� /      Meeting     P|	�/V  �}	�/V  �m	Some_stuffs_Some_stuffs_ /V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  Xs��$�K� /      Appointment `'	�/V  �(	�/V  �)	This_stuffs_This_stuffs_ /V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  �R	�/V  T	�/V  p����
�W� /       Workout     P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ���-� �lٳ /      Some_stuffs p��/V  ���/V  ��This_stuffs_This_stuffs_ /V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �/V  P�/V  ���-� ��۳ /      Birthday    ��/V  p�/V  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  ���-� ��ڳ /      Some_stuffs Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  Q ��cw1K� /      Some_stuffs  �ҿ&V  p�ҿ&V  0��justforfun_justforfun_ ҿ&V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  R ��cw1��� /      Some_stuffs P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  S ��cw1K� /      Some_stuffs  U�/V  pW�/V  0Yjustforfun_justforfun_ �/V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  !�u�m.d~
 /      Workout     ���/V   ��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  ��(~�m.��
 /      Some_stuffs � �/V  0�/V  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  p�K�n.n /      Meeting /V  p��/V  ���/V  ��This_stuffs_This_stuffs_ /V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  �5U�n._) /      Meeting     P$�/V  �%�/V   'This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  (|��n.�S /       Appointment PIӿ&V  �Jӿ&V  �M�Some_stuffs_Some_stuffs_ &V  �Vӿ&V  @Xӿ&V  p[ӿ&V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  9�_��n.g� /       Birthday    ��/V  p�/V  pjustforfun_justforfun_ �/V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  ���Ko._ /      Workout     ���/V  ���/V   �Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V   ����o.$� /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �1���o.p' /      Birthday V  � �/V  0�/V  pjustforfun_justforfun_ �/V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  q���p."R /      Birthday    �e�/V  �f�/V  0]Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  8��(\x.'� /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �~�Ēx.� /      Workout     P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �:�x.�� /   	   Some_stuffs ���/V   ��/V  ��Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �/V  P�/V  ��/V  �/V  ��׬�y.� /      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �-�Дz.�' /      Meeting     ���/V   ��/V  `�This_stuffs_This_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  ��u9Ƃ.q�* /       Meeting                        justforfun_justforfun_                                                                                                                                                                                                                                               �4���.��* /      Birthday                       This_stuffs_This_stuffs_                                                                                                                                                                                                                                             I��x�.Ù+ /      Meeting     ���/V  ���/V  @�justforfun_justforfun_ 	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  ��Sv��.v�+ /      Workout                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     @ؔ\��.(^, /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �vb�1�.��, /       Meeting /V  0s�/V  pt�/V  �uThis_stuffs_This_stuffs_ /V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  �����.�G- /      Meeting     P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ����+�.��8 /      Meeting     P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  	�����.��9 /      Meeting /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  C&L�.�: /      Birthday V   U�/V  pW�/V  0Yjustforfun_justforfun_ �/V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �؉tE�.�f: /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     a�7���.�u; /      Some_stuffs P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �)��.w�; /      Meeting /V  ���/V   ��/V  `�justforfun_justforfun_ �/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  �Ƽ^a�.�< /      Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     k����.�^< /      Birthday    ��/V  `�/V  �#Some_stuffs_Some_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  ������.��H /      Workout     PIӿ&V  �Jӿ&V  �M�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �K�<)�.YI /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �1mw�.:�I /      Appointment  U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  a�2\ݗ.LiJ /      Birthday    P�/V  PQ�/V  0HThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  �C�%y�.�TK /       Appointment  U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  9�U&�.G�V /      Birthday V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  iҠ�A�.�W /      Meeting     0s�/V  pt�/V  �uThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  q��H\�.N@W /      Appointment �Z�/V  �[�/V  �RSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V  Hk�	��.ɯW /       Workout     �	�/V  �/V  PSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �,����.�Y /      Workout     �#�/V  P%�/V  �)This_stuffs_This_stuffs_ /V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V   =����.`�Y /      Appointment                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     x��'H�.�'Z /      Appointment `FԿ&V  �GԿ&V  `I�This_stuffs_This_stuffs_ &V  �NԿ&V  �VԿ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  @      E!]�.cGZ /      Appointment ���/V  ���/V  p�This_stuffs_This_stuffs_ /V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �\���.��Z /       Birthday V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  ��:Ţ.��Z /      Some_stuffs � �/V  0�/V  pThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  ��/?�.Q1f /      Some_stuffs �z�/V  ���/V  �~Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  �0�iq�.>}f /      Workout /V  �	�/V  �/V  PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �r���.>�f /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               @�E��.Hhg /       Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     x0U�>�.��g /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               `��Z��.��h /      Meeting     PIӿ&V  �Jӿ&V  �M�Some_stuffs_Some_stuffs_ &V  �Vӿ&V  @Xӿ&V  p[ӿ&V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �`>�.�uj /       Workout     P�/V  PQ�/V  0Hjustforfun_justforfun_ �/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  Yl�椴.\�u /      Birthday    0]�/V  p^�/V  �_This_stuffs_This_stuffs_ /V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  �Pش.�5v /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �{ς?�.��v /      Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             X�%N��.�Hw /      Meeting     ���/V  @��/V  p�Some_stuffs_Some_stuffs_ /V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  ��µ.��w /      Appointment P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��_7��.X�w /      Some_stuffs  <�/V  �F�/V  @?Some_stuffs_Some_stuffs_ /V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  �A��.Bx /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ���x�.�x /      Birthday    ���/V  @��/V  p�This_stuffs_This_stuffs_ /V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  1^{�:�.Fd� /      Workout /V  ���/V  0��/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  @      �+���.5�� /      Meeting /V  � �/V  0�/V  pThis_stuffs_This_stuffs_ /V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  ��Ȇ>�.6� /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               +i��.�� /   	   Workout     P�/V  PQ�/V  0HSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  (���.�_� /       Appointment ���/V   ��/V  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V  h�@
��.m�� /   	   Birthday    �ӿ&V  `�ӿ&V  ���This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  @�ӿ&V  ��ӿ&V  p�ӿ&V  0�ӿ&V  p�ӿ&V  @�ӿ&V  ��ӿ&V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  ��g��.�i� /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               �x#V�.�-� /      Appointment ��/V  p�/V  pThis_stuffs_This_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  Q��ܾ�.*̕ /      Meeting     ��/V   �/V  p+This_stuffs_This_stuffs_ /V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  .I�W�.㲖 /      Meeting     м�/V  ��/V  @�This_stuffs_This_stuffs_ /V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  �N����.� /   	   Appointment  ��/V  @��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���4��.�W� /       Meeting /V  P 
�/V  �
�/V  
This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  
�/V  �$
�/V  �%
�/V   
�/V  `
�/V  �
�/V  
�/V  P
�/V  �
�/V  P
�/V  �
�/V  �
�/V  
�/V  P
�/V  � 
�/V  "
�/V  :
�/V   '
�/V  `(
�/V  �)
�/V  �*
�/V   ,
�/V  �-
�/V   /
�/V  `0
�/V  �1
�/V  Q�Kt@�.�� /      Workout     ��/V  `�/V  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  ��[�.:;� /      Birthday V  0~Կ&V  pԿ&V  �x�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  `�Կ&V  ��Կ&V  @�Կ&V  @�Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  ��Կ&V  `�Կ&V  ��Կ&V  `�Կ&V  0�Կ&V  p�Կ&V   �Կ&V  @�Կ&V  ��Կ&V   �Կ&V  P�Կ&V  ��Կ&V  �Կ&V  0�Կ&V  p�Կ&V  �Կ&V  `�Կ&V  ���`��.8>� /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ��,8��.��� /      Workout     ���/V   ��/V  `�This_stuffs_This_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  1W�@&�.f�� /      Appointment ���/V   ��/V  `�This_stuffs_This_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  @�.���.�|� /      Some_stuffs PIӿ&V  �Jӿ&V  �M�justforfun_justforfun_ ӿ&V  �Vӿ&V  @Xӿ&V  p[ӿ&V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �$G���.ݵ� /       Appointment  �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  A9��"�.�� /      Workout     `��/V  ���/V  0�justforfun_justforfun_ �/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  �-T=�.CŴ /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             Y�q���.K�� /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ���%�.�$� /      Meeting     �Z�/V  �[�/V  �RSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V  q��;p�6 ȥ /       Birthday V  �	�/V  P	�/V  �		This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  r��;p�6 9� /      Some_stuffs                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             s��;p�6 �� /   	   Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     t��;p�6 � /   	   Appointment  �ҿ&V  p�ҿ&V  0��justforfun_justforfun_ ҿ&V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  u��;p�6 ȥ /       Birthday    PIӿ&V  �Jӿ&V  �M�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ &V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  v��;p�6 9� /      Some_stuffs ��/V  p�/V  pThis_stuffs_This_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  w��;p�6 �� /   	   Workout     ���/V  ���/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  @+`���%�z� /       Some_stuffs ���/V  @��/V  p�Some_stuffs_Some_stuffs_ /V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  (���t�#.�� /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               q����#.� /       Birthday    Ј�/V  P��/V  ЏThis_stuffs_This_stuffs_ /V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  r����#.) /   	   Appointment ���/V  ���/V  �Some_stuffs_Some_stuffs_ /V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  )�U��#.�O /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             *�U��#.�S /       Appointment @��/V  ���/V  ��Some_stuffs_Some_stuffs_ /V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @      !��m$.5� /   	   Some_stuffs ���/V  ���/V   �This_stuffs_This_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  "��m$.$� /      Birthday V  P�/V  ��/V  justforfun_justforfun_ �/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �c1�w$.�* /      Birthday V  PZ	�/V  �[	�/V  `L	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �c1�w$.�& /      Birthday    `�/V  ��/V  �	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �R>�N�$.3p /      Appointment P$�/V  �%�/V   'justforfun_justforfun_ �/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  9>�^�'.�� /      Meeting     � �/V  0�/V  pjustforfun_justforfun_ �/V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V  :>�^�'.�� /      Birthday    ��	�/V  0�	�/V  p�	Some_stuffs_Some_stuffs_ /V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  �
�/V  �
�/V  ��	�/V  �	�/V  P 
�/V  �
�/V  
�/V  P
�/V  �
�/V  
�/V  �
�/V  

�/V  �
�/V  
�/V  �$
�/V  �%
�/V   
�/V  `
�/V  �
�/V  
�/V  P
�/V  �
�/V  P
�/V  �r�'�(.�. /      Appointment �	�/V  0�	�/V  p�	Some_stuffs_Some_stuffs_ /V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  p�	�/V  @�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  �c�@K(.�� /      Workout     ��/V  p�/V  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  �c�@K(.� /      Workout      ��/V  @��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ��8��+.��* /      Appointment  U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ��8��+.q�* /       Meeting     P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ���/�+.M+ /      Birthday    �	�/V  0�	�/V  p�	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  0�	�/V  p�	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  p�	�/V  @�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ��	�/V  ��	�/V  0�	�/V  p�	�/V  ���/�+.� + /      Workout     ��/V  0��/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  �qW�),.��+ /      Birthday    P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  �qW�),.v�+ /      Workout      ��/V  @��/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  AEtשF,.�[, /      Birthday    Ј�/V  P��/V  ЏThis_stuffs_This_stuffs_ /V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  BEtשF,.(^, /      Some_stuffs  U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ����,.�B- /      Some_stuffs ���/V  ���/V   �Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  ����,.rK- /      Birthday     ��/V  `��/V  мSome_stuffs_Some_stuffs_ /V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  `k�.t�/.l9 /      Appointment ���/V  P��/V  �Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V  ���i7�/.�c: /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             ���i7�/.�f: /      Appointment �	�/V  �/V  PSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  ��:�B0.��; /      Some_stuffs �
�/V  
�/V  P
Some_stuffs_Some_stuffs_ /V   '
�/V  `(
�/V  �)
�/V  �*
�/V   ,
�/V  �-
�/V   /
�/V  `0
�/V  �1
�/V  `3
�/V  �4
�/V   6
�/V  �7
�/V  �N
�/V  P;
�/V  �<
�/V  >
�/V  �?
�/V  A
�/V  PB
�/V  �C
�/V  �D
�/V  F
�/V  PG
�/V  �H
�/V  �I
�/V  K
�/V  �L
�/V  �c
�/V  ��j�V0.E< /       Workout /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ��j�V0.�< /      Workout     P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ���Ej3.��G /      Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ��K���3.��H /      Some_stuffs Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  ��K���3.��H /      Workout     ���/V   ��/V  @�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ���/V   ��/V  `��/V  0��/V  p��/V  ���/V  �-F:��3.<�H /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             ����1�3.J_I /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ����1�3.YI /      Birthday V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �z%�hG4.�SK /       Workout     �$	�/V   &	�/V  `'	Some_stuffs_Some_stuffs_ /V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  07	�/V  �8	�/V   K	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  �z%�hG4.�XK /   	   Meeting     ���/V  Ъ�/V  P�justforfun_justforfun_ �/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V  0�~��e4.��K /      Meeting     0H�/V  pI�/V  �JSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  I�8�x7.d�W /      Appointment P$�/V  �%�/V   'This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  J�8�x7.Y�W /       Appointment @@	�/V  �A	�/V  �B	justforfun_justforfun_ 	�/V  �G	�/V  0I	�/V  PZ	�/V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  h��>h�7.�X /      Appointment `��/V  ���/V  0�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  �/y��7.\�X /      Some_stuffs ��/V  P��/V  ��justforfun_justforfun_ �/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  �n��7.��X /      Meeting                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �T��3�7.�Y /   	   Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               �T��3�7. Y /      Workout                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �@q-�7.��Y /      Appointment �z�/V  ���/V  �~justforfun_justforfun_ �/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  �@q-�7.`�Y /      Appointment ���/V  P��/V  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V  yz�E8.>&Z /      Workout     �	�/V  �/V  PThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  zz�E8.�'Z /      Appointment ��/V   �/V  �!This_stuffs_This_stuffs_ /V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  PQ�/V  0H�/V  �}Gw$8.�HZ /      Appointment �#�/V  P%�/V  �)This_stuffs_This_stuffs_ /V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  �}Gw$8.MZ /      Workout                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ��eێ98._�Z /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ��eێ98.��Z /       Birthday V  ��/V  P��/V  ��This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  p���V8.�	[ /   	   Some_stuffs ��/V  p�/V  pThis_stuffs_This_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  �%F��.;.�	f /      Some_stuffs  U�/V  pW�/V  0Yjustforfun_justforfun_ �/V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �����8;./f /      Meeting     0s�/V  pt�/V  �uThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  �����8;.�1f /      Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �'�]b;.\�f /      Workout     ��	�/V  П	�/V  `�	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  P�	�/V  ��	�/V  Л	�/V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  Ю	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  �'�]b;. �f /      Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  A@o$�;.�lg /      Workout /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  B@o$�;.Hhg /       Meeting /V   <�/V  �F�/V  @?Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  y�\���;.ɳg /      Workout     ��/V  p�/V  pSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  z�\���;.��g /      Appointment ���/V  0��/V  p�justforfun_justforfun_ �/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  0/E*i�;.&xh /      Meeting     P|	�/V  �}	�/V  �m	This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V  ��	�/V  П	�/V  `�	�/V  ��	�/V  �	�/V  P�	�/V  ��	�/V  Ж	�/V  �	�/V  P�	�/V  ��	�/V  aP!��;.�h /       Some_stuffs `M�/V  �N�/V  �ZThis_stuffs_This_stuffs_ /V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  bP!��;.��h /      Meeting /V  @��/V  ���/V  ��Some_stuffs_Some_stuffs_ /V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �J�P�;.��h /      Meeting     P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/��?.o�v /       Workout     Ј�/V  P��/V  ЏThis_stuffs_This_stuffs_ /V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  ��/��?.��v /      Appointment ���/V  0��/V  p�Some_stuffs_Some_stuffs_ /V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  ���/V   ��/V  `��/V  м�/V  Y?�X��?.EEw /      Appointment @@	�/V  �A	�/V  �B	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  Z?�X��?.,Kw /   	   Appointment  U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V   �
��?.�x /      Workout /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V   �
��?.Bx /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �9<B�?.�x /      Birthday    ��/V  p�/V  pSome_stuffs_Some_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  �9<B�?.�x /      Workout     ���/V  @��/V  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  ����lC.u� /   	   Workout /V  �	�/V  �/V  PSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   �/V  �!�/V  #�/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  ����lC.6� /      Birthday     ��/V  @��/V  ��justforfun_justforfun_ �/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  ipkD.�� /      Workout     ���/V  @��/V  p�Some_stuffs_Some_stuffs_ /V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ��/V  ��/V  `�/V  @�/V  ��/V  ��/V  jpkD.m�� /   	   Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     ����G.qՓ /      Appointment P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ���+G.�m� /      Some_stuffs  U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  ���+G.�i� /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               �å�'H.p=� /      Birthday    ���/V  ���/V  p�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �å�'H.:;� /      Birthday V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �3�f�K.:�� /      Meeting     �		�/V  �
	�/V  	justforfun_justforfun_ 	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  �Ǜ��;K.%� /      Meeting     P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ���#OK.=o� /      Appointment 0]�/V  p^�/V  �_Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  ���/V  �~�/V   ��/V  @��/V  ���/V  ���/V  0��/V  p��/V  P��/V  ���/V  0��/V  p��/V  �)q�mK.� /      Birthday    ���/V   ��/V  @�This_stuffs_This_stuffs_ /V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  �	�/V  `	�/V  �	�/V  �	�/V  P	�/V  �		�/V  �
	�/V  	�/V  P	�/V  �	�/V  p	�/V  �	�/V   	�/V  `	�/V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V  A�}_�N.Kx� /      Birthday    ��/V  `�/V  �#This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  B�}_�N.�|� /      Some_stuffs ��/V  `�/V  �justforfun_justforfun_ �/V  ��/V  `�/V  ��/V   �/V  p+�/V  �,�/V  P$�/V  �%�/V   '�/V  @(�/V  �)�/V  @5�/V  �-�/V  p/�/V  �0�/V  p2�/V  �3�/V   >�/V  �6�/V   8�/V  �9�/V  �:�/V   <�/V  �F�/V  @?�/V  �@�/V  @B�/V  �C�/V  P�/V  ���u�AO.{�� /   	   Workout     p��/V  ���/V  ��Some_stuffs_Some_stuffs_ /V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �/V  P�/V  ���u�AO.ݵ� /       Appointment ���/V  P��/V  �This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  @��/V  ���/V  ���/V  ���/V  ��/V  P��/V  ���/V  ���/V  ��/V  P��/V  ���/V   ��/V  ���/V  0��/V  p��/V  ���/V   ��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V  ��O�IKO.0ڳ /      Some_stuffs                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     ���O.�Ǵ /      Birthday    P��/V  Ъ�/V  ЭSome_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  ���O.CŴ /      Some_stuffs ���/V   ��/V  `�Some_stuffs_Some_stuffs_ /V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  P�����O.J�� /   	   Meeting     Ј�/V  P��/V  ЏSome_stuffs_Some_stuffs_ /V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  �E���S0�"� /       Meeting /V   U�/V  pW�/V  0YThis_stuffs_This_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  �{K�T9dx� /      Appointment Ј�/V  P��/V  Џjustforfun_justforfun_ �/V   ��/V  @��/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  �{K�T9�r� /      Meeting     ���/V  ���/V  p�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �{K�T9#q� /      Birthday                       This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �{K�T9dx� /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               AW�;n3GE�� /      Workout                        justforfun_justforfun_                                                                                                                                                                                                                                               BW�;n3G�� /       Appointment ��/V  p�/V  pSome_stuffs_Some_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  CW�;n3GE�� /      Workout     `M�/V  �N�/V  �Zjustforfun_justforfun_ �/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  �v�/V  0x�/V  py�/V  �z�/V  DW�;n3G)�� /   	   Some_stuffs `��/V  ���/V  `�This_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  p��/V   ��/V  @��/V  ���/V   ��/V  P�/V  ��/V  � �/V  0�/V  p�/V  ��/V  `�/V  ��/V  �	�/V  �/V  P�/V  ��/V  �/V  ��/V  ��/V  `�/V  ��/V   �/V  �!�/V  #�/V  ��/V  EW�;n3G��� /      Meeting     �		�/V  �
	�/V  	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �	�/V  	�/V  P	�/V  �	�/V  �	�/V  @	�/V  �,	�/V  �	�/V   !	�/V  `"	�/V  �#	�/V  �$	�/V   &	�/V  `'	�/V  �(	�/V  �)	�/V  P+	�/V  ;	�/V  P<	�/V  �-	�/V  @/	�/V  �0	�/V   2	�/V  @3	�/V  �4	�/V  �5	�/V  I�"�XƄYW� /      Workout      ��/V  @��/V  ��Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  @��/V  ���/V  `��/V  ��/V  `��/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  ���/V   ��/V  ���/V   ��/V  @��/V  ���/V   ��/V   ��/V  ���/V   ��/V  @��/V  @��/V  ���/V  @��/V  ���/V  ���/V  J�"�XƄYR� /      Meeting     ��/V  `�/V  �#Some_stuffs_Some_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  K�"�XƄY�� /      Some_stuffs ��ӿ&V  p�ӿ&V  0��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  L�"�XƄYW� /      Workout &V  PIӿ&V  �Jӿ&V  �M�Some_stuffs_Some_stuffs_ &V  �Vӿ&V  @Xӿ&V  p[ӿ&V  �\ӿ&V  0`ӿ&V  �aӿ&V   eӿ&V  �fӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  qt�Z�Ha /      Workout     ��/V  p�/V  pThis_stuffs_This_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  rt�Z�Ha߽� /   	   Birthday V  ��
�/V  ��
�/V  0�
This_stuffs_This_stuffs_ /V  ��
�/V   �
�/V  `�
�/V  ��
�/V  ��
�/V   �
�/V  P�
�/V  ��
�/V  Е
�/V  P�
�/V  ��
�/V  Й
�/V  �
�/V  ��
�/V  �
�/V  ��
�/V  Р
�/V  �
�/V  p�
�/V  ��
�/V  �
�/V  0�
�/V  @�
�/V  ��
�/V  @�
�/V  ��
�/V   �
�/V  @�
�/V  ��
�/V  st�Z�Ha��� /      Birthday                       Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             tt�Z�HaN�� /       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     p�����k� /      Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             y.唕�$l� /      Workout      ��/V  ���/V  ��justforfun_justforfun_ �/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V   ��/V  ���/V  ���/V  @��/V  � 	�/V  �	�/V  z.唕�$l� /      Appointment ���/V  0��/V  p�Some_stuffs_Some_stuffs_ /V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  0��/V  p��/V  {.唕�$l� /      Meeting &V   �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  |.唕�$l/� /   	   Some_stuffs p[ӿ&V  �\ӿ&V  0`�Some_stuffs_Some_stuffs_ &V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  Y�p�'�v�� /      Meeting /V  �Q	�/V  �R	�/V  T	Some_stuffs_Some_stuffs_ /V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  Z�p�'�vF� /      Birthday    P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  [�p�'�v�� /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               \�p�'�vK� /      Appointment ��ӿ&V  p�ӿ&V  0��This_stuffs_This_stuffs_ &V  `�ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  ��ӿ&V  P�ӿ&V  `Կ&V  �Կ&V  �Կ&V  @	Կ&V  pԿ&V  �Կ&V  0Կ&V  pԿ&V  �Կ&V  �Կ&V   "Կ&V  `#Կ&V  �(Կ&V  P*Կ&V  �/Կ&V  P1Կ&V  �6Կ&V  `8Կ&V   >Կ&V  @?Կ&V  �9Կ&V   ;Կ&V  �<Կ&V  �a�N�dx�� /      Appointment �/�/V   1�/V  �5Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  P��/V  ���/V  `��/V   ��/V  	�7��f��"+ /      Meeting      <�/V  �F�/V  @?justforfun_justforfun_ �/V  P�/V  PQ�/V  0H�/V  pI�/V  �J�/V   L�/V  `M�/V  �N�/V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V  
�7��f�$+ /      Workout     �0	�/V   2	�/V  @3	Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �7��f�%+ /   	   Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             �7��f�a#+ /      Meeting                        Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             i�L�����ow /      Some_stuffs ��/V  p�/V  pSome_stuffs_Some_stuffs_ /V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  j�L�����nw /   	   Some_stuffs ��/V  p�/V  pjustforfun_justforfun_ �/V  ��/V  `�/V  �#�/V  P%�/V  �)�/V  P+�/V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  k�L����-mw /       Some_stuffs                    This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     l�L�����ow /      Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             A��cg˥�8�w /      Appointment P��/V  Ъ�/V  Эjustforfun_justforfun_ �/V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  B��cg˥�,�w /      Workout /V   U�/V  pW�/V  0YSome_stuffs_Some_stuffs_ /V   b�/V  �c�/V  �f�/V   h�/V  k�/V  �l�/V  �n�/V   p�/V  @r�/V  �t�/V  x�/V  �y�/V  �{�/V  P}�/V  ��/V   ��/V  ���/V  ���/V  ���/V  p��/V   ��/V  ���/V  ��/V  ���/V  @��/V  ���/V  p��/V  ��/V  ���/V  C��cg˥�C�w /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               D��cg˥���w /      Appointment                    Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     �Z�����+ /      Workout     @3	�/V  �4	�/V  �5	justforfun_justforfun_ 	�/V  �=	�/V  �>	�/V  @@	�/V  �A	�/V  �B	�/V  0D	�/V  pE	�/V  �F	�/V  �G	�/V  0I	�/V  PZ	�/V  �[	�/V  `L	�/V  �M	�/V  �N	�/V   P	�/V  �Q	�/V  �R	�/V  T	�/V  PU	�/V  �V	�/V   X	�/V   k	�/V  `l	�/V  �\	�/V  ^	�/V  �_	�/V  �`	�/V  `b	�/V  �Z����ͼ+ /      Meeting     ��	�/V  Ж	�/V  �	Some_stuffs_Some_stuffs_ /V  �	�/V  P�	�/V  �	�/V  0�	�/V  �	�/V  P�	�/V  ��	�/V  Ф	�/V  �	�/V  P�	�/V  ��	�/V  Щ	�/V  �	�/V  P�	�/V  ��	�/V  Ю	�/V  ��	�/V   �	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  0�	�/V  p�	�/V  ��	�/V  �	�/V  �Z����"�+ /      Appointment                    This_stuffs_This_stuffs_                                                                                                                                                                                                                                             �Z����"�+ /   	   Meeting                        Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     AM8��g+�Pz� /      Workout     P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_ /V  ���/V  @��/V  p��/V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  BM8��g+��x� /      Birthday                       justforfun_justforfun_                                                                                                                                                                                                                                               CM8��g+�/}� /   	   Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             DM8��g+��z� /       Some_stuffs                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             EM8��g+�Pz� /      Workout                        This_stuffs_This_stuffs_                                                                                                                                                                                                                                             !��������r- /      Some_stuffs ��/V  `�/V  �#Some_stuffs_Some_stuffs_ /V  �/�/V   1�/V  �5�/V  @7�/V  �;�/V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  "�������Wq- /      Meeting     p��/V  P��/V  ��This_stuffs_This_stuffs_ /V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  ���/V  Ю�/V  ��/V  ���/V  P��/V  ��/V  #��������r- /      Appointment                    justforfun_justforfun_                                                                                                                                                                                                                                               $��������r- /      Some_stuffs  �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �E��fa���(� /      Some_stuffs ���/V   ��/V  ��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V   ��/V  ���/V  ���/V  @��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V  0��/V  ���/V  ���/V  ��/V  ���/V  ���/V   ��/V  @��/V  ���/V  ���/V   ��/V  @��/V   	�/V  0��/V  ���/V  ���/V  �E��fa���(� /      Meeting                        This_stuffs_This_stuffs_This_stuffs_This_stuffs_                                                                                                                                                                                                                     �E��fa���"� /       Meeting &V   �ҿ&V  p�ҿ&V  0��This_stuffs_This_stuffs_ &V   ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �E��fa���(� /      Some_stuffs  �ҿ&V  p�ҿ&V  0��Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ &V   ӿ&V  ӿ&V  �ӿ&V  �ӿ&V   ӿ&V  @ӿ&V  �ӿ&V  ӿ&V  �ӿ&V  �ӿ&V  Pӿ&V  �ӿ&V   !ӿ&V  �#ӿ&V  �$ӿ&V  �&ӿ&V  p(ӿ&V   ,ӿ&V  �-ӿ&V  0ӿ&V  �2ӿ&V  @5ӿ&V  �6ӿ&V  p9ӿ&V  �:ӿ&V  �=ӿ&V  �E��fa�Ǡ+� /      Some_stuffs ���/V  ���/V   �Some_stuffs_Some_stuffs_ /V  ���/V   ��/V  `��/V  ���/V  0��/V  p��/V  ���/V  ���/V  p��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ���/V  @��/V  @��/V  ���/V  `��/V  ���/V  `��/V  ���/V  ���/V  `��/V  ���/V  `��/V  0��/V  p��/V   ��/V  �E��fa���(� /      Meeting     P��/V  Ъ�/V  ЭThis_stuffs_This_stuffs_This_stuffs_This_stuffs_ /V  ��/V  0��/V  ���/V   ��/V  ���/V  ���/V  `��/V  ���/V  ���/V  P��/V  ���/V  `��/V  ���/V  @��/V  ���/V  p��/V  ���/V  0��/V  ���/V  ���/V   ��/V  ���/V  `��/V  ��/V  ���/V  ���/V  @�o2$:��裗 /      Appointment �~�/V   ��/V  @�Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  0��/V  p��/V  ���/V  ���/V  0��/V  p��/V  0��/V  ���/V  Д�/V  ��/V  P��/V  ���/V  Й�/V  ��/V  P��/V  p��/V  ���/V  ��/V  p��/V  ��/V   ��/V  `��/V  ���/V  ���/V  Ъ�/V  P��/V  q�-��q��X� /      Birthday    �#�/V  P%�/V  �)Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_ /V  p=�/V  0B�/V  pC�/V  @H�/V  �I�/V  `N�/V  �O�/V  �T�/V  V�/V  �Z�/V  P\�/V  `a�/V  �b�/V  �g�/V  @i�/V  pn�/V  �o�/V  0u�/V  pv�/V  �{�/V  �|�/V   ��/V  `��/V  Ј�/V  P��/V  Џ�/V  r�-��q�*X� /      Workout     0H�/V  pI�/V  �JSome_stuffs_Some_stuffs_ /V  �Z�/V  �[�/V  �R�/V  �S�/V  U�/V  PV�/V  �W�/V  �X�/V  �e�/V  �f�/V  0]�/V  p^�/V  �_�/V  �`�/V  0b�/V  pc�/V  �p�/V  �q�/V  h�/V  �i�/V  �j�/V   l�/V  @m�/V  �n�/V  |�/V  P}�/V  0s�/V  pt�/V  �u�/V  s�-��q�GT� /      Birthday                       Some_stuffs_Some_stuffs_Some_stuffs_Some_stuffs_                                                                                                                                                                                                                     t�-��q�W� /       Workout &V  `IԿ&V  �PԿ&V   L�justforfun_justforfun_ Կ&V   RԿ&V  �SԿ&V   UԿ&V  �\Կ&V   XԿ&V  @YԿ&V  �ZԿ&V   cԿ&V   ^Կ&V  �_Կ&V   aԿ&V  @iԿ&V  @dԿ&V  �eԿ&V  @gԿ&V  �oԿ&V  �jԿ&V  �kԿ&V   mԿ&V  `nԿ&V  0vԿ&V  pwԿ&V  �pԿ&V   rԿ&V  `sԿ&V  �tԿ&V  0~Կ&V  pԿ&V  �xԿ&V  A�����%�x�f /   	   Some_stuffs  k	�/V  `l	�/V  �\	Some_stuffs_Some_stuffs_ /V  `b	�/V  �c	�/V  e	�/V  Pf	�/V  �g	�/V  �h	�/V  P|	�/V  �}	�/V  �m	�/V  �n	�/V  Pp	�/V  �q	�/V   s	�/V  @t	�/V  �u	�/V  �v	�/V  `x	�/V  �y	�/V  ��	�/V   �	�/V  �~	�/V  @�	�/V  ��	�/V  ��	�/V   �	�/V  @�	�/V  ��	�/V   �	�/V  @�	�/V  B�����%��f /      Birthday     �	�/V  `�	�/V  ��	justforfun_justforfun_ 	�/V  p�	�/V  ��	�/V  0�	�/V  ��	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  ��	�/V  0�	�/V  �
�/V  �
�/V  ��	�/V  �	�/V  P 
�/V  �
�/V  
�/V  P
�/V  �
�/V  
�/V  �
�/V  

�/V  �
�/V  
�/V  �$
�/V  �%
�/V   
�/V  `
�/V  �
�/V  C�����%f /       Appointment                    Some_stuffs_Some_stuffs_                                                                                                                                                                                                                                             D�����%�ȣf /      Appointment p[ӿ&V  �\ӿ&V  0`�justforfun_justforfun_ ӿ&V  �iӿ&V  `kӿ&V  �nӿ&V  �oӿ&V  Psӿ&V  �tӿ&V  `xӿ&V  �yӿ&V  @}ӿ&V  �~ӿ&V  p�ӿ&V  ��ӿ&V  0�ӿ&V  ��ӿ&V  ��ӿ&V   �ӿ&V  ��ӿ&V  `�ӿ&V  �ӿ&V  ��ӿ&V  ��ӿ&V  �ӿ&V  �ӿ&V  `�ӿ&V  @�ӿ&V  ��ӿ&V  �ӿ&V  p�ӿ&V  p�ӿ&V  